// Chris Ceroici 

module RNE(
	S0, S1, S2, S3, S4, S5, S6, S7, S8, S9, S10, S11, S12, S13, S14, S15, S16, S17, S18, S19, S20, S21, S22, S23, S24, S25, S26, S27, S28, S29, S30, S31, S32, S33, S34, S35, S36, S37, S38, S39, S40, S41, S42, S43, S44, S45, S46, S47, S48, S49, S50, S51, S52, S53, S54, S55, S56, S57, S58, S59, S60, S61, S62, S63, S64, S65, S66, S67, S68, S69, S70, S71, S72, S73, S74, S75, S76, S77, S78, S79, S80, S81, S82, S83, S84, S85, S86, S87, S88, S89, S90, S91, S92, S93, S94, S95, S96, S97, S98, S99, S100, S101, S102, S103, S104, S105, S106, S107, S108, S109, S110, S111, S112, S113, S114, S115, S116, S117, S118, S119, S120, S121, S122, S123, S124, S125, S126, S127, S128, S129, S130, S131, S132, S133, S134, S135, S136, S137, S138, S139, S140, S141, S142, S143, S144, S145, S146, S147, S148, S149, S150, S151, S152, S153, S154, S155, S156, S157, S158, S159, S160, S161, S162, S163, S164, S165, S166, S167, S168, S169, S170, S171, S172, S173, S174, S175, S176, S177, S178, S179, S180, S181, S182, S183, S184, S185, S186, S187, S188, S189, S190, S191, S192, S193, S194, S195, S196, S197, S198, S199, S200, S201, S202, S203, S204, S205, S206, S207, S208, S209, S210, S211, S212, S213, S214, S215, S216, S217, S218, S219, S220, S221, S222, S223, S224, S225, S226, S227, S228, S229, S230, S231, S232, S233, S234, S235, S236, S237, S238, S239, S240, S241, S242, S243, S244, S245, S246, S247, S248, S249, S250, S251, S252, S253, S254, S255, S256, S257, S258, S259, S260, S261, S262, S263, S264, S265, S266, S267, S268, S269, S270, S271, S272, S273, S274, S275, S276, S277, S278, S279,
	R0, R1, R2, R3, R4, R5, R6, R7, R8, R9, R10, R11, R12, R13, R14, R15, R16, R17, R18, R19, R20, R21, R22, R23, R24, R25, R26, R27, R28, R29, R30, R31, R32, R33, R34, R35, R36, R37, R38, R39, R40, R41, R42, R43, R44, R45, R46, R47, R48, R49, R50, R51, R52, R53, R54, R55, R56, R57, R58, R59, R60, R61, R62, R63, R64, R65, R66, R67, R68, R69, R70, R71, R72, R73, R74, R75, R76, R77, R78, R79, R80, R81, R82, R83, R84, R85, R86, R87, R88, R89, R90, R91, R92, R93, R94, R95, R96, R97, R98, R99, R100, R101, R102, R103, R104, R105, R106, R107, R108, R109, R110, R111, R112, R113, R114, R115, R116, R117, R118, R119, R120, R121, R122, R123, R124, R125, R126, R127, R128, R129, R130, R131, R132, R133, R134, R135, R136, R137, R138, R139, R140, R141, R142, R143, R144, R145, R146, R147, R148, R149, R150, R151, R152, R153, R154, R155, R156, R157, R158, R159, R160, R161, R162, R163, R164, R165, R166, R167, R168, R169, R170, R171, R172, R173, R174, R175, R176, R177, R178, R179, R180, R181, R182, R183, R184, R185, R186, R187, R188, R189, R190, R191, R192, R193, R194, R195, R196, R197, R198, R199, R200, R201, R202, R203, R204, R205, R206, R207, R208, R209, R210, R211, R212, R213, R214, R215, R216, R217, R218, R219, R220, R221, R222, R223, R224, R225, R226, R227, R228, R229, R230, R231, R232, R233, R234, R235, R236, R237, R238, R239, R240, R241, R242, R243, R244, R245, R246, R247, R248, R249, R250, R251, R252, R253, R254, R255, R256, R257, R258, R259, R260, R261, R262, R263, R264, R265, R266, R267, R268, R269, R270, R271, R272, R273, R274, R275, R276, R277, R278, R279, R280, R281, R282, R283, R284, R285, R286, R287, R288, R289, R290, R291, R292, R293, R294, R295, R296, R297, R298, R299, R300, R301, R302, R303, R304, R305, R306, R307, R308, R309, R310, R311, R312, R313, R314, R315, R316, R317, R318, R319, R320, R321, R322, R323, R324, R325, R326, R327, R328, R329, R330, R331, R332, R333, R334, R335, R336, R337, R338, R339, R340, R341, R342, R343, R344, R345, R346, R347, R348, R349, R350, R351, R352, R353, R354, R355, R356, R357, R358, R359, R360, R361, R362, R363, R364, R365, R366, R367, R368, R369, R370, R371, R372, R373, R374, R375, R376, R377, R378, R379, R380, R381, R382, R383, R384, R385, R386, R387, R388, R389, R390, R391, R392, R393, R394, R395, R396, R397, R398, R399, R400, R401, R402, R403, R404, R405, R406, R407, R408, R409, R410, R411, R412, R413, R414, R415, R416, R417, R418, R419, R420, R421, R422, R423, R424, R425, R426, R427, R428, R429, R430, R431, R432, R433, R434, R435, R436, R437, R438, R439, R440, R441, R442, R443, R444, R445, R446, R447, R448, R449, R450, R451, R452, R453, R454, R455, R456, R457, R458, R459, R460, R461, R462, R463, R464, R465, R466, R467, R468, R469, R470, R471, R472, R473, R474, R475, R476, R477, R478, R479, R480, R481, R482, R483, R484, R485, R486, R487, R488, R489, R490, R491, R492, R493, R494, R495, R496, R497, R498, R499, R500, R501, R502, R503, R504, R505, R506, R507, R508, R509, R510, R511, R512, R513, R514, R515, R516, R517, R518, R519, R520, R521, R522, R523, R524, R525, R526, R527, R528,
	R_long0, R_long1, R_long2, R_long3, R_long4, R_long5, R_long6, R_long7, R_long8, R_long9, R_long10, R_long11, R_long12, R_long13, R_long14,
	CLK, INIT_powerup, SDcount
); 

parameter DP = 8; // RN precision
parameter DPlong =16; // RN alpha precision
parameter LFSR_S = 16; // LFSR size

input CLK, INIT_powerup; // Initialization signal (new set)
input [31:0] SDcount;
input wire [16 - 1:0] S0, S1, S2, S3, S4, S5, S6, S7, S8, S9, S10, S11, S12, S13, S14, S15, S16, S17, S18, S19, S20, S21, S22, S23, S24, S25, S26, S27, S28, S29, S30, S31, S32, S33, S34, S35, S36, S37, S38, S39, S40, S41, S42, S43, S44, S45, S46, S47, S48, S49, S50, S51, S52, S53, S54, S55, S56, S57, S58, S59, S60, S61, S62, S63, S64, S65, S66, S67, S68, S69, S70, S71, S72, S73, S74, S75, S76, S77, S78, S79, S80, S81, S82, S83, S84, S85, S86, S87, S88, S89, S90, S91, S92, S93, S94, S95, S96, S97, S98, S99, S100, S101, S102, S103, S104, S105, S106, S107, S108, S109, S110, S111, S112, S113, S114, S115, S116, S117, S118, S119, S120, S121, S122, S123, S124, S125, S126, S127, S128, S129, S130, S131, S132, S133, S134, S135, S136, S137, S138, S139, S140, S141, S142, S143, S144, S145, S146, S147, S148, S149, S150, S151, S152, S153, S154, S155, S156, S157, S158, S159, S160, S161, S162, S163, S164, S165, S166, S167, S168, S169, S170, S171, S172, S173, S174, S175, S176, S177, S178, S179, S180, S181, S182, S183, S184, S185, S186, S187, S188, S189, S190, S191, S192, S193, S194, S195, S196, S197, S198, S199, S200, S201, S202, S203, S204, S205, S206, S207, S208, S209, S210, S211, S212, S213, S214, S215, S216, S217, S218, S219, S220, S221, S222, S223, S224, S225, S226, S227, S228, S229, S230, S231, S232, S233, S234, S235, S236, S237, S238, S239, S240, S241, S242, S243, S244, S245, S246, S247, S248, S249, S250, S251, S252, S253, S254, S255, S256, S257, S258, S259, S260, S261, S262, S263, S264, S265, S266, S267, S268, S269, S270, S271, S272, S273, S274, S275, S276, S277, S278, S279;
output [DP - 1:0] R0, R1, R2, R3, R4, R5, R6, R7, R8, R9, R10, R11, R12, R13, R14, R15, R16, R17, R18, R19, R20, R21, R22, R23, R24, R25, R26, R27, R28, R29, R30, R31, R32, R33, R34, R35, R36, R37, R38, R39, R40, R41, R42, R43, R44, R45, R46, R47, R48, R49, R50, R51, R52, R53, R54, R55, R56, R57, R58, R59, R60, R61, R62, R63, R64, R65, R66, R67, R68, R69, R70, R71, R72, R73, R74, R75, R76, R77, R78, R79, R80, R81, R82, R83, R84, R85, R86, R87, R88, R89, R90, R91, R92, R93, R94, R95, R96, R97, R98, R99, R100, R101, R102, R103, R104, R105, R106, R107, R108, R109, R110, R111, R112, R113, R114, R115, R116, R117, R118, R119, R120, R121, R122, R123, R124, R125, R126, R127, R128, R129, R130, R131, R132, R133, R134, R135, R136, R137, R138, R139, R140, R141, R142, R143, R144, R145, R146, R147, R148, R149, R150, R151, R152, R153, R154, R155, R156, R157, R158, R159, R160, R161, R162, R163, R164, R165, R166, R167, R168, R169, R170, R171, R172, R173, R174, R175, R176, R177, R178, R179, R180, R181, R182, R183, R184, R185, R186, R187, R188, R189, R190, R191, R192, R193, R194, R195, R196, R197, R198, R199, R200, R201, R202, R203, R204, R205, R206, R207, R208, R209, R210, R211, R212, R213, R214, R215, R216, R217, R218, R219, R220, R221, R222, R223, R224, R225, R226, R227, R228, R229, R230, R231, R232, R233, R234, R235, R236, R237, R238, R239, R240, R241, R242, R243, R244, R245, R246, R247, R248, R249, R250, R251, R252, R253, R254, R255, R256, R257, R258, R259, R260, R261, R262, R263, R264, R265, R266, R267, R268, R269, R270, R271, R272, R273, R274, R275, R276, R277, R278, R279, R280, R281, R282, R283, R284, R285, R286, R287, R288, R289, R290, R291, R292, R293, R294, R295, R296, R297, R298, R299, R300, R301, R302, R303, R304, R305, R306, R307, R308, R309, R310, R311, R312, R313, R314, R315, R316, R317, R318, R319, R320, R321, R322, R323, R324, R325, R326, R327, R328, R329, R330, R331, R332, R333, R334, R335, R336, R337, R338, R339, R340, R341, R342, R343, R344, R345, R346, R347, R348, R349, R350, R351, R352, R353, R354, R355, R356, R357, R358, R359, R360, R361, R362, R363, R364, R365, R366, R367, R368, R369, R370, R371, R372, R373, R374, R375, R376, R377, R378, R379, R380, R381, R382, R383, R384, R385, R386, R387, R388, R389, R390, R391, R392, R393, R394, R395, R396, R397, R398, R399, R400, R401, R402, R403, R404, R405, R406, R407, R408, R409, R410, R411, R412, R413, R414, R415, R416, R417, R418, R419, R420, R421, R422, R423, R424, R425, R426, R427, R428, R429, R430, R431, R432, R433, R434, R435, R436, R437, R438, R439, R440, R441, R442, R443, R444, R445, R446, R447, R448, R449, R450, R451, R452, R453, R454, R455, R456, R457, R458, R459, R460, R461, R462, R463, R464, R465, R466, R467, R468, R469, R470, R471, R472, R473, R474, R475, R476, R477, R478, R479, R480, R481, R482, R483, R484, R485, R486, R487, R488, R489, R490, R491, R492, R493, R494, R495, R496, R497, R498, R499, R500, R501, R502, R503, R504, R505, R506, R507, R508, R509, R510, R511, R512, R513, R514, R515, R516, R517, R518, R519, R520, R521, R522, R523, R524, R525, R526, R527, R528;
output [DPlong - 1:0] R_long0, R_long1, R_long2, R_long3, R_long4, R_long5, R_long6, R_long7, R_long8, R_long9, R_long10, R_long11, R_long12, R_long13, R_long14;

wire [DP-1:0] R529,R530,R531,R532,R533,R534,R535,R536,R537,R538,R539,R540,R541,R542,R543;

// Short RN LFSRs
cascLFSR_16Tap xLFSR0(.TRIG(CLK),.RESET(INIT_powerup),.OUT0(R0),.OUT1(R527),.OUT2(R32),.OUT3(R495),.OUT4(R64),.OUT5(R463),.OUT6(R96),.OUT7(R431),.OUT8(R128),.OUT9(R399),.OUT10(R160),.OUT11(R367),.OUT12(R192),.OUT13(R335),.OUT14(R224),.OUT15(R303),.SEED(S0), .SDcount(SDcount)); 
cascLFSR_16Tap xLFSR1(.TRIG(CLK),.RESET(INIT_powerup),.OUT0(R256),.OUT1(R271),.OUT2(R288),.OUT3(R239),.OUT4(R320),.OUT5(R207),.OUT6(R352),.OUT7(R175),.OUT8(R384),.OUT9(R143),.OUT10(R416),.OUT11(R111),.OUT12(R448),.OUT13(R79),.OUT14(R480),.OUT15(R47),.SEED(S8), .SDcount(SDcount)); 
cascLFSR_16Tap xLFSR2(.TRIG(CLK),.RESET(INIT_powerup),.OUT0(R512),.OUT1(R15),.OUT2(R1),.OUT3(R526),.OUT4(R33),.OUT5(R494),.OUT6(R65),.OUT7(R462),.OUT8(R97),.OUT9(R430),.OUT10(R129),.OUT11(R398),.OUT12(R161),.OUT13(R366),.OUT14(R193),.OUT15(R334),.SEED(S16), .SDcount(SDcount)); 
cascLFSR_16Tap xLFSR3(.TRIG(CLK),.RESET(INIT_powerup),.OUT0(R225),.OUT1(R302),.OUT2(R257),.OUT3(R270),.OUT4(R289),.OUT5(R238),.OUT6(R321),.OUT7(R206),.OUT8(R353),.OUT9(R174),.OUT10(R385),.OUT11(R142),.OUT12(R417),.OUT13(R110),.OUT14(R449),.OUT15(R78),.SEED(S24), .SDcount(SDcount)); 
cascLFSR_16Tap xLFSR4(.TRIG(CLK),.RESET(INIT_powerup),.OUT0(R481),.OUT1(R46),.OUT2(R513),.OUT3(R14),.OUT4(R2),.OUT5(R525),.OUT6(R34),.OUT7(R493),.OUT8(R66),.OUT9(R461),.OUT10(R98),.OUT11(R429),.OUT12(R130),.OUT13(R397),.OUT14(R162),.OUT15(R365),.SEED(S32), .SDcount(SDcount)); 
cascLFSR_16Tap xLFSR5(.TRIG(CLK),.RESET(INIT_powerup),.OUT0(R194),.OUT1(R333),.OUT2(R226),.OUT3(R301),.OUT4(R258),.OUT5(R269),.OUT6(R290),.OUT7(R237),.OUT8(R322),.OUT9(R205),.OUT10(R354),.OUT11(R173),.OUT12(R386),.OUT13(R141),.OUT14(R418),.OUT15(R109),.SEED(S40), .SDcount(SDcount)); 
cascLFSR_16Tap xLFSR6(.TRIG(CLK),.RESET(INIT_powerup),.OUT0(R450),.OUT1(R77),.OUT2(R482),.OUT3(R45),.OUT4(R514),.OUT5(R13),.OUT6(R3),.OUT7(R524),.OUT8(R35),.OUT9(R492),.OUT10(R67),.OUT11(R460),.OUT12(R99),.OUT13(R428),.OUT14(R131),.OUT15(R396),.SEED(S48), .SDcount(SDcount)); 
cascLFSR_16Tap xLFSR7(.TRIG(CLK),.RESET(INIT_powerup),.OUT0(R163),.OUT1(R364),.OUT2(R195),.OUT3(R332),.OUT4(R227),.OUT5(R300),.OUT6(R259),.OUT7(R268),.OUT8(R291),.OUT9(R236),.OUT10(R323),.OUT11(R204),.OUT12(R355),.OUT13(R172),.OUT14(R387),.OUT15(R140),.SEED(S56), .SDcount(SDcount)); 
cascLFSR_16Tap xLFSR8(.TRIG(CLK),.RESET(INIT_powerup),.OUT0(R419),.OUT1(R108),.OUT2(R451),.OUT3(R76),.OUT4(R483),.OUT5(R44),.OUT6(R515),.OUT7(R12),.OUT8(R4),.OUT9(R523),.OUT10(R36),.OUT11(R491),.OUT12(R68),.OUT13(R459),.OUT14(R100),.OUT15(R427),.SEED(S64), .SDcount(SDcount)); 
cascLFSR_16Tap xLFSR9(.TRIG(CLK),.RESET(INIT_powerup),.OUT0(R132),.OUT1(R395),.OUT2(R164),.OUT3(R363),.OUT4(R196),.OUT5(R331),.OUT6(R228),.OUT7(R299),.OUT8(R260),.OUT9(R267),.OUT10(R292),.OUT11(R235),.OUT12(R324),.OUT13(R203),.OUT14(R356),.OUT15(R171),.SEED(S72), .SDcount(SDcount)); 
cascLFSR_16Tap xLFSR10(.TRIG(CLK),.RESET(INIT_powerup),.OUT0(R388),.OUT1(R139),.OUT2(R420),.OUT3(R107),.OUT4(R452),.OUT5(R75),.OUT6(R484),.OUT7(R43),.OUT8(R516),.OUT9(R11),.OUT10(R5),.OUT11(R522),.OUT12(R37),.OUT13(R490),.OUT14(R69),.OUT15(R458),.SEED(S80), .SDcount(SDcount)); 
cascLFSR_16Tap xLFSR11(.TRIG(CLK),.RESET(INIT_powerup),.OUT0(R101),.OUT1(R426),.OUT2(R133),.OUT3(R394),.OUT4(R165),.OUT5(R362),.OUT6(R197),.OUT7(R330),.OUT8(R229),.OUT9(R298),.OUT10(R261),.OUT11(R266),.OUT12(R293),.OUT13(R234),.OUT14(R325),.OUT15(R202),.SEED(S88), .SDcount(SDcount)); 
cascLFSR_16Tap xLFSR12(.TRIG(CLK),.RESET(INIT_powerup),.OUT0(R357),.OUT1(R170),.OUT2(R389),.OUT3(R138),.OUT4(R421),.OUT5(R106),.OUT6(R453),.OUT7(R74),.OUT8(R485),.OUT9(R42),.OUT10(R517),.OUT11(R10),.OUT12(R6),.OUT13(R521),.OUT14(R38),.OUT15(R489),.SEED(S96), .SDcount(SDcount)); 
cascLFSR_16Tap xLFSR13(.TRIG(CLK),.RESET(INIT_powerup),.OUT0(R70),.OUT1(R457),.OUT2(R102),.OUT3(R425),.OUT4(R134),.OUT5(R393),.OUT6(R166),.OUT7(R361),.OUT8(R198),.OUT9(R329),.OUT10(R230),.OUT11(R297),.OUT12(R262),.OUT13(R265),.OUT14(R294),.OUT15(R233),.SEED(S104), .SDcount(SDcount)); 
cascLFSR_16Tap xLFSR14(.TRIG(CLK),.RESET(INIT_powerup),.OUT0(R326),.OUT1(R201),.OUT2(R358),.OUT3(R169),.OUT4(R390),.OUT5(R137),.OUT6(R422),.OUT7(R105),.OUT8(R454),.OUT9(R73),.OUT10(R486),.OUT11(R41),.OUT12(R518),.OUT13(R9),.OUT14(R7),.OUT15(R520),.SEED(S112), .SDcount(SDcount)); 
cascLFSR_16Tap xLFSR15(.TRIG(CLK),.RESET(INIT_powerup),.OUT0(R39),.OUT1(R488),.OUT2(R71),.OUT3(R456),.OUT4(R103),.OUT5(R424),.OUT6(R135),.OUT7(R392),.OUT8(R167),.OUT9(R360),.OUT10(R199),.OUT11(R328),.OUT12(R231),.OUT13(R296),.OUT14(R263),.OUT15(R264),.SEED(S120), .SDcount(SDcount)); 
cascLFSR_16Tap xLFSR16(.TRIG(CLK),.RESET(INIT_powerup),.OUT0(R295),.OUT1(R232),.OUT2(R327),.OUT3(R200),.OUT4(R359),.OUT5(R168),.OUT6(R391),.OUT7(R136),.OUT8(R423),.OUT9(R104),.OUT10(R455),.OUT11(R72),.OUT12(R487),.OUT13(R40),.OUT14(R519),.OUT15(R8),.SEED(S128), .SDcount(SDcount)); 
cascLFSR_16Tap xLFSR17(.TRIG(CLK),.RESET(INIT_powerup),.OUT0(R535),.OUT1(R24),.OUT2(R503),.OUT3(R56),.OUT4(R471),.OUT5(R88),.OUT6(R439),.OUT7(R120),.OUT8(R407),.OUT9(R152),.OUT10(R375),.OUT11(R184),.OUT12(R343),.OUT13(R216),.OUT14(R311),.OUT15(R248),.SEED(S136), .SDcount(SDcount)); 
cascLFSR_16Tap xLFSR18(.TRIG(CLK),.RESET(INIT_powerup),.OUT0(R279),.OUT1(R280),.OUT2(R247),.OUT3(R312),.OUT4(R215),.OUT5(R344),.OUT6(R183),.OUT7(R376),.OUT8(R151),.OUT9(R408),.OUT10(R119),.OUT11(R440),.OUT12(R87),.OUT13(R472),.OUT14(R55),.OUT15(R504),.SEED(S144), .SDcount(SDcount)); 
cascLFSR_16Tap xLFSR19(.TRIG(CLK),.RESET(INIT_powerup),.OUT0(R23),.OUT1(R536),.OUT2(R534),.OUT3(R25),.OUT4(R502),.OUT5(R57),.OUT6(R470),.OUT7(R89),.OUT8(R438),.OUT9(R121),.OUT10(R406),.OUT11(R153),.OUT12(R374),.OUT13(R185),.OUT14(R342),.OUT15(R217),.SEED(S152), .SDcount(SDcount)); 
cascLFSR_16Tap xLFSR20(.TRIG(CLK),.RESET(INIT_powerup),.OUT0(R310),.OUT1(R249),.OUT2(R278),.OUT3(R281),.OUT4(R246),.OUT5(R313),.OUT6(R214),.OUT7(R345),.OUT8(R182),.OUT9(R377),.OUT10(R150),.OUT11(R409),.OUT12(R118),.OUT13(R441),.OUT14(R86),.OUT15(R473),.SEED(S160), .SDcount(SDcount)); 
cascLFSR_16Tap xLFSR21(.TRIG(CLK),.RESET(INIT_powerup),.OUT0(R54),.OUT1(R505),.OUT2(R22),.OUT3(R537),.OUT4(R533),.OUT5(R26),.OUT6(R501),.OUT7(R58),.OUT8(R469),.OUT9(R90),.OUT10(R437),.OUT11(R122),.OUT12(R405),.OUT13(R154),.OUT14(R373),.OUT15(R186),.SEED(S168), .SDcount(SDcount)); 
cascLFSR_16Tap xLFSR22(.TRIG(CLK),.RESET(INIT_powerup),.OUT0(R341),.OUT1(R218),.OUT2(R309),.OUT3(R250),.OUT4(R277),.OUT5(R282),.OUT6(R245),.OUT7(R314),.OUT8(R213),.OUT9(R346),.OUT10(R181),.OUT11(R378),.OUT12(R149),.OUT13(R410),.OUT14(R117),.OUT15(R442),.SEED(S176), .SDcount(SDcount)); 
cascLFSR_16Tap xLFSR23(.TRIG(CLK),.RESET(INIT_powerup),.OUT0(R85),.OUT1(R474),.OUT2(R53),.OUT3(R506),.OUT4(R21),.OUT5(R538),.OUT6(R532),.OUT7(R27),.OUT8(R500),.OUT9(R59),.OUT10(R468),.OUT11(R91),.OUT12(R436),.OUT13(R123),.OUT14(R404),.OUT15(R155),.SEED(S184), .SDcount(SDcount)); 
cascLFSR_16Tap xLFSR24(.TRIG(CLK),.RESET(INIT_powerup),.OUT0(R372),.OUT1(R187),.OUT2(R340),.OUT3(R219),.OUT4(R308),.OUT5(R251),.OUT6(R276),.OUT7(R283),.OUT8(R244),.OUT9(R315),.OUT10(R212),.OUT11(R347),.OUT12(R180),.OUT13(R379),.OUT14(R148),.OUT15(R411),.SEED(S192), .SDcount(SDcount)); 
cascLFSR_16Tap xLFSR25(.TRIG(CLK),.RESET(INIT_powerup),.OUT0(R116),.OUT1(R443),.OUT2(R84),.OUT3(R475),.OUT4(R52),.OUT5(R507),.OUT6(R20),.OUT7(R539),.OUT8(R531),.OUT9(R28),.OUT10(R499),.OUT11(R60),.OUT12(R467),.OUT13(R92),.OUT14(R435),.OUT15(R124),.SEED(S200), .SDcount(SDcount)); 
cascLFSR_16Tap xLFSR26(.TRIG(CLK),.RESET(INIT_powerup),.OUT0(R403),.OUT1(R156),.OUT2(R371),.OUT3(R188),.OUT4(R339),.OUT5(R220),.OUT6(R307),.OUT7(R252),.OUT8(R275),.OUT9(R284),.OUT10(R243),.OUT11(R316),.OUT12(R211),.OUT13(R348),.OUT14(R179),.OUT15(R380),.SEED(S208), .SDcount(SDcount)); 
cascLFSR_16Tap xLFSR27(.TRIG(CLK),.RESET(INIT_powerup),.OUT0(R147),.OUT1(R412),.OUT2(R115),.OUT3(R444),.OUT4(R83),.OUT5(R476),.OUT6(R51),.OUT7(R508),.OUT8(R19),.OUT9(R540),.OUT10(R530),.OUT11(R29),.OUT12(R498),.OUT13(R61),.OUT14(R466),.OUT15(R93),.SEED(S216), .SDcount(SDcount)); 
cascLFSR_16Tap xLFSR28(.TRIG(CLK),.RESET(INIT_powerup),.OUT0(R434),.OUT1(R125),.OUT2(R402),.OUT3(R157),.OUT4(R370),.OUT5(R189),.OUT6(R338),.OUT7(R221),.OUT8(R306),.OUT9(R253),.OUT10(R274),.OUT11(R285),.OUT12(R242),.OUT13(R317),.OUT14(R210),.OUT15(R349),.SEED(S224), .SDcount(SDcount)); 
cascLFSR_16Tap xLFSR29(.TRIG(CLK),.RESET(INIT_powerup),.OUT0(R178),.OUT1(R381),.OUT2(R146),.OUT3(R413),.OUT4(R114),.OUT5(R445),.OUT6(R82),.OUT7(R477),.OUT8(R50),.OUT9(R509),.OUT10(R18),.OUT11(R541),.OUT12(R529),.OUT13(R30),.OUT14(R497),.OUT15(R62),.SEED(S232), .SDcount(SDcount)); 
cascLFSR_16Tap xLFSR30(.TRIG(CLK),.RESET(INIT_powerup),.OUT0(R465),.OUT1(R94),.OUT2(R433),.OUT3(R126),.OUT4(R401),.OUT5(R158),.OUT6(R369),.OUT7(R190),.OUT8(R337),.OUT9(R222),.OUT10(R305),.OUT11(R254),.OUT12(R273),.OUT13(R286),.OUT14(R241),.OUT15(R318),.SEED(S240), .SDcount(SDcount)); 
cascLFSR_16Tap xLFSR31(.TRIG(CLK),.RESET(INIT_powerup),.OUT0(R209),.OUT1(R350),.OUT2(R177),.OUT3(R382),.OUT4(R145),.OUT5(R414),.OUT6(R113),.OUT7(R446),.OUT8(R81),.OUT9(R478),.OUT10(R49),.OUT11(R510),.OUT12(R17),.OUT13(R542),.OUT14(R528),.OUT15(R31),.SEED(S248), .SDcount(SDcount)); 
cascLFSR_16Tap xLFSR32(.TRIG(CLK),.RESET(INIT_powerup),.OUT0(R496),.OUT1(R63),.OUT2(R464),.OUT3(R95),.OUT4(R432),.OUT5(R127),.OUT6(R400),.OUT7(R159),.OUT8(R368),.OUT9(R191),.OUT10(R336),.OUT11(R223),.OUT12(R304),.OUT13(R255),.OUT14(R272),.OUT15(R287),.SEED(S256), .SDcount(SDcount)); 
cascLFSR_16Tap xLFSR33(.TRIG(CLK),.RESET(INIT_powerup),.OUT0(R240),.OUT1(R319),.OUT2(R208),.OUT3(R351),.OUT4(R176),.OUT5(R383),.OUT6(R144),.OUT7(R415),.OUT8(R112),.OUT9(R447),.OUT10(R80),.OUT11(R479),.OUT12(R48),.OUT13(R511),.OUT14(R16),.OUT15(R543),.SEED(S264), .SDcount(SDcount)); 

// Long RN LFSRs
cascLFSR xLFSR_L0(.TRIG(CLK),.RESET(INIT_powerup),.OUT1(R_long0[7:0]),.OUT2(R_long0[15:8]),.SEED(S265),.SDcount(SDcount));
cascLFSR xLFSR_L1(.TRIG(CLK),.RESET(INIT_powerup),.OUT1(R_long1[7:0]),.OUT2(R_long1[15:8]),.SEED(S266),.SDcount(SDcount));
cascLFSR xLFSR_L2(.TRIG(CLK),.RESET(INIT_powerup),.OUT1(R_long2[7:0]),.OUT2(R_long2[15:8]),.SEED(S267),.SDcount(SDcount));
cascLFSR xLFSR_L3(.TRIG(CLK),.RESET(INIT_powerup),.OUT1(R_long3[7:0]),.OUT2(R_long3[15:8]),.SEED(S268),.SDcount(SDcount));
cascLFSR xLFSR_L4(.TRIG(CLK),.RESET(INIT_powerup),.OUT1(R_long4[7:0]),.OUT2(R_long4[15:8]),.SEED(S269),.SDcount(SDcount));
cascLFSR xLFSR_L5(.TRIG(CLK),.RESET(INIT_powerup),.OUT1(R_long5[7:0]),.OUT2(R_long5[15:8]),.SEED(S270),.SDcount(SDcount));
cascLFSR xLFSR_L6(.TRIG(CLK),.RESET(INIT_powerup),.OUT1(R_long6[7:0]),.OUT2(R_long6[15:8]),.SEED(S271),.SDcount(SDcount));
cascLFSR xLFSR_L7(.TRIG(CLK),.RESET(INIT_powerup),.OUT1(R_long7[7:0]),.OUT2(R_long7[15:8]),.SEED(S272),.SDcount(SDcount));
cascLFSR xLFSR_L8(.TRIG(CLK),.RESET(INIT_powerup),.OUT1(R_long8[7:0]),.OUT2(R_long8[15:8]),.SEED(S273),.SDcount(SDcount));
cascLFSR xLFSR_L9(.TRIG(CLK),.RESET(INIT_powerup),.OUT1(R_long9[7:0]),.OUT2(R_long9[15:8]),.SEED(S274),.SDcount(SDcount));
cascLFSR xLFSR_L10(.TRIG(CLK),.RESET(INIT_powerup),.OUT1(R_long10[7:0]),.OUT2(R_long10[15:8]),.SEED(S275),.SDcount(SDcount));
cascLFSR xLFSR_L11(.TRIG(CLK),.RESET(INIT_powerup),.OUT1(R_long11[7:0]),.OUT2(R_long11[15:8]),.SEED(S276),.SDcount(SDcount));
cascLFSR xLFSR_L12(.TRIG(CLK),.RESET(INIT_powerup),.OUT1(R_long12[7:0]),.OUT2(R_long12[15:8]),.SEED(S277),.SDcount(SDcount));
cascLFSR xLFSR_L13(.TRIG(CLK),.RESET(INIT_powerup),.OUT1(R_long13[7:0]),.OUT2(R_long13[15:8]),.SEED(S278),.SDcount(SDcount));
cascLFSR xLFSR_L14(.TRIG(CLK),.RESET(INIT_powerup),.OUT1(R_long14[7:0]),.OUT2(R_long14[15:8]),.SEED(S279),.SDcount(SDcount));

endmodule
