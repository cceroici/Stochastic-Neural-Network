// Chris Ceroici

// Parallel network training evaluator
// Version 9.0

module NETPAR_GRADIENT(
	dalpha_L1_j_0_netPar0, dalpha_L1_j_1_netPar0, dalpha_L1_j_2_netPar0, dalpha_L1_j_3_netPar0, dalpha_L1_j_4_netPar0, dalpha_L1_j_5_netPar0, dalpha_L1_j_6_netPar0, dalpha_L1_j_7_netPar0, dalpha_L1_j_8_netPar0, dalpha_L1_j_9_netPar0, dalpha_L1_j_10_netPar0, dalpha_L1_j_11_netPar0, dalpha_L1_j_12_netPar0, dalpha_L1_j_13_netPar0, dalpha_L1_j_14_netPar0, dalpha_L1_j_15_netPar0, dalpha_L1_j_16_netPar0, dalpha_L1_j_17_netPar0, dalpha_L1_j_18_netPar0, dalpha_L1_j_19_netPar0, dalpha_L1_j_20_netPar0, dalpha_L1_j_21_netPar0, dalpha_L1_j_22_netPar0, dalpha_L1_j_23_netPar0, dalpha_L1_j_24_netPar0,
	dbeta_L1_netPar0,
	dalpha_L2_j_0_netPar0, dalpha_L2_j_1_netPar0, dalpha_L2_j_2_netPar0, dalpha_L2_j_3_netPar0, dalpha_L2_j_4_netPar0, dalpha_L2_j_5_netPar0, dalpha_L2_j_6_netPar0, dalpha_L2_j_7_netPar0,
	dbeta_L2_netPar0,
	dalpha_L3_j_0_netPar0, dalpha_L3_j_1_netPar0, dalpha_L3_j_2_netPar0, dalpha_L3_j_3_netPar0, dalpha_L3_j_4_netPar0,
	dbeta_L3_netPar0,
	SIGN_dalpha_L1_j_0_netPar0, SIGN_dalpha_L1_j_1_netPar0, SIGN_dalpha_L1_j_2_netPar0, SIGN_dalpha_L1_j_3_netPar0, SIGN_dalpha_L1_j_4_netPar0, SIGN_dalpha_L1_j_5_netPar0, SIGN_dalpha_L1_j_6_netPar0, SIGN_dalpha_L1_j_7_netPar0, SIGN_dalpha_L1_j_8_netPar0, SIGN_dalpha_L1_j_9_netPar0, SIGN_dalpha_L1_j_10_netPar0, SIGN_dalpha_L1_j_11_netPar0, SIGN_dalpha_L1_j_12_netPar0, SIGN_dalpha_L1_j_13_netPar0, SIGN_dalpha_L1_j_14_netPar0, SIGN_dalpha_L1_j_15_netPar0, SIGN_dalpha_L1_j_16_netPar0, SIGN_dalpha_L1_j_17_netPar0, SIGN_dalpha_L1_j_18_netPar0, SIGN_dalpha_L1_j_19_netPar0, SIGN_dalpha_L1_j_20_netPar0, SIGN_dalpha_L1_j_21_netPar0, SIGN_dalpha_L1_j_22_netPar0, SIGN_dalpha_L1_j_23_netPar0, SIGN_dalpha_L1_j_24_netPar0,
	SIGN_dbeta_L1_netPar0,
	SIGN_dalpha_L2_j_0_netPar0, SIGN_dalpha_L2_j_1_netPar0, SIGN_dalpha_L2_j_2_netPar0, SIGN_dalpha_L2_j_3_netPar0, SIGN_dalpha_L2_j_4_netPar0, SIGN_dalpha_L2_j_5_netPar0, SIGN_dalpha_L2_j_6_netPar0, SIGN_dalpha_L2_j_7_netPar0,
	SIGN_dbeta_L2_netPar0,
	SIGN_dalpha_L3_j_0_netPar0, SIGN_dalpha_L3_j_1_netPar0, SIGN_dalpha_L3_j_2_netPar0, SIGN_dalpha_L3_j_3_netPar0, SIGN_dalpha_L3_j_4_netPar0,
	SIGN_dbeta_L3_netPar0,
	dalpha_L1_j_0_netPar1, dalpha_L1_j_1_netPar1, dalpha_L1_j_2_netPar1, dalpha_L1_j_3_netPar1, dalpha_L1_j_4_netPar1, dalpha_L1_j_5_netPar1, dalpha_L1_j_6_netPar1, dalpha_L1_j_7_netPar1, dalpha_L1_j_8_netPar1, dalpha_L1_j_9_netPar1, dalpha_L1_j_10_netPar1, dalpha_L1_j_11_netPar1, dalpha_L1_j_12_netPar1, dalpha_L1_j_13_netPar1, dalpha_L1_j_14_netPar1, dalpha_L1_j_15_netPar1, dalpha_L1_j_16_netPar1, dalpha_L1_j_17_netPar1, dalpha_L1_j_18_netPar1, dalpha_L1_j_19_netPar1, dalpha_L1_j_20_netPar1, dalpha_L1_j_21_netPar1, dalpha_L1_j_22_netPar1, dalpha_L1_j_23_netPar1, dalpha_L1_j_24_netPar1,
	dbeta_L1_netPar1,
	dalpha_L2_j_0_netPar1, dalpha_L2_j_1_netPar1, dalpha_L2_j_2_netPar1, dalpha_L2_j_3_netPar1, dalpha_L2_j_4_netPar1, dalpha_L2_j_5_netPar1, dalpha_L2_j_6_netPar1, dalpha_L2_j_7_netPar1,
	dbeta_L2_netPar1,
	dalpha_L3_j_0_netPar1, dalpha_L3_j_1_netPar1, dalpha_L3_j_2_netPar1, dalpha_L3_j_3_netPar1, dalpha_L3_j_4_netPar1,
	dbeta_L3_netPar1,
	SIGN_dalpha_L1_j_0_netPar1, SIGN_dalpha_L1_j_1_netPar1, SIGN_dalpha_L1_j_2_netPar1, SIGN_dalpha_L1_j_3_netPar1, SIGN_dalpha_L1_j_4_netPar1, SIGN_dalpha_L1_j_5_netPar1, SIGN_dalpha_L1_j_6_netPar1, SIGN_dalpha_L1_j_7_netPar1, SIGN_dalpha_L1_j_8_netPar1, SIGN_dalpha_L1_j_9_netPar1, SIGN_dalpha_L1_j_10_netPar1, SIGN_dalpha_L1_j_11_netPar1, SIGN_dalpha_L1_j_12_netPar1, SIGN_dalpha_L1_j_13_netPar1, SIGN_dalpha_L1_j_14_netPar1, SIGN_dalpha_L1_j_15_netPar1, SIGN_dalpha_L1_j_16_netPar1, SIGN_dalpha_L1_j_17_netPar1, SIGN_dalpha_L1_j_18_netPar1, SIGN_dalpha_L1_j_19_netPar1, SIGN_dalpha_L1_j_20_netPar1, SIGN_dalpha_L1_j_21_netPar1, SIGN_dalpha_L1_j_22_netPar1, SIGN_dalpha_L1_j_23_netPar1, SIGN_dalpha_L1_j_24_netPar1,
	SIGN_dbeta_L1_netPar1,
	SIGN_dalpha_L2_j_0_netPar1, SIGN_dalpha_L2_j_1_netPar1, SIGN_dalpha_L2_j_2_netPar1, SIGN_dalpha_L2_j_3_netPar1, SIGN_dalpha_L2_j_4_netPar1, SIGN_dalpha_L2_j_5_netPar1, SIGN_dalpha_L2_j_6_netPar1, SIGN_dalpha_L2_j_7_netPar1,
	SIGN_dbeta_L2_netPar1,
	SIGN_dalpha_L3_j_0_netPar1, SIGN_dalpha_L3_j_1_netPar1, SIGN_dalpha_L3_j_2_netPar1, SIGN_dalpha_L3_j_3_netPar1, SIGN_dalpha_L3_j_4_netPar1,
	SIGN_dbeta_L3_netPar1,
	dalpha_L1_j_0_netPar2, dalpha_L1_j_1_netPar2, dalpha_L1_j_2_netPar2, dalpha_L1_j_3_netPar2, dalpha_L1_j_4_netPar2, dalpha_L1_j_5_netPar2, dalpha_L1_j_6_netPar2, dalpha_L1_j_7_netPar2, dalpha_L1_j_8_netPar2, dalpha_L1_j_9_netPar2, dalpha_L1_j_10_netPar2, dalpha_L1_j_11_netPar2, dalpha_L1_j_12_netPar2, dalpha_L1_j_13_netPar2, dalpha_L1_j_14_netPar2, dalpha_L1_j_15_netPar2, dalpha_L1_j_16_netPar2, dalpha_L1_j_17_netPar2, dalpha_L1_j_18_netPar2, dalpha_L1_j_19_netPar2, dalpha_L1_j_20_netPar2, dalpha_L1_j_21_netPar2, dalpha_L1_j_22_netPar2, dalpha_L1_j_23_netPar2, dalpha_L1_j_24_netPar2,
	dbeta_L1_netPar2,
	dalpha_L2_j_0_netPar2, dalpha_L2_j_1_netPar2, dalpha_L2_j_2_netPar2, dalpha_L2_j_3_netPar2, dalpha_L2_j_4_netPar2, dalpha_L2_j_5_netPar2, dalpha_L2_j_6_netPar2, dalpha_L2_j_7_netPar2,
	dbeta_L2_netPar2,
	dalpha_L3_j_0_netPar2, dalpha_L3_j_1_netPar2, dalpha_L3_j_2_netPar2, dalpha_L3_j_3_netPar2, dalpha_L3_j_4_netPar2,
	dbeta_L3_netPar2,
	SIGN_dalpha_L1_j_0_netPar2, SIGN_dalpha_L1_j_1_netPar2, SIGN_dalpha_L1_j_2_netPar2, SIGN_dalpha_L1_j_3_netPar2, SIGN_dalpha_L1_j_4_netPar2, SIGN_dalpha_L1_j_5_netPar2, SIGN_dalpha_L1_j_6_netPar2, SIGN_dalpha_L1_j_7_netPar2, SIGN_dalpha_L1_j_8_netPar2, SIGN_dalpha_L1_j_9_netPar2, SIGN_dalpha_L1_j_10_netPar2, SIGN_dalpha_L1_j_11_netPar2, SIGN_dalpha_L1_j_12_netPar2, SIGN_dalpha_L1_j_13_netPar2, SIGN_dalpha_L1_j_14_netPar2, SIGN_dalpha_L1_j_15_netPar2, SIGN_dalpha_L1_j_16_netPar2, SIGN_dalpha_L1_j_17_netPar2, SIGN_dalpha_L1_j_18_netPar2, SIGN_dalpha_L1_j_19_netPar2, SIGN_dalpha_L1_j_20_netPar2, SIGN_dalpha_L1_j_21_netPar2, SIGN_dalpha_L1_j_22_netPar2, SIGN_dalpha_L1_j_23_netPar2, SIGN_dalpha_L1_j_24_netPar2,
	SIGN_dbeta_L1_netPar2,
	SIGN_dalpha_L2_j_0_netPar2, SIGN_dalpha_L2_j_1_netPar2, SIGN_dalpha_L2_j_2_netPar2, SIGN_dalpha_L2_j_3_netPar2, SIGN_dalpha_L2_j_4_netPar2, SIGN_dalpha_L2_j_5_netPar2, SIGN_dalpha_L2_j_6_netPar2, SIGN_dalpha_L2_j_7_netPar2,
	SIGN_dbeta_L2_netPar2,
	SIGN_dalpha_L3_j_0_netPar2, SIGN_dalpha_L3_j_1_netPar2, SIGN_dalpha_L3_j_2_netPar2, SIGN_dalpha_L3_j_3_netPar2, SIGN_dalpha_L3_j_4_netPar2,
	SIGN_dbeta_L3_netPar2,
	dalpha_L1_j_0, dalpha_L1_j_1, dalpha_L1_j_2, dalpha_L1_j_3, dalpha_L1_j_4, dalpha_L1_j_5, dalpha_L1_j_6, dalpha_L1_j_7, dalpha_L1_j_8, dalpha_L1_j_9, dalpha_L1_j_10, dalpha_L1_j_11, dalpha_L1_j_12, dalpha_L1_j_13, dalpha_L1_j_14, dalpha_L1_j_15, dalpha_L1_j_16, dalpha_L1_j_17, dalpha_L1_j_18, dalpha_L1_j_19, dalpha_L1_j_20, dalpha_L1_j_21, dalpha_L1_j_22, dalpha_L1_j_23, dalpha_L1_j_24,
	dbeta_L1,
	dalpha_L2_j_0, dalpha_L2_j_1, dalpha_L2_j_2, dalpha_L2_j_3, dalpha_L2_j_4, dalpha_L2_j_5, dalpha_L2_j_6, dalpha_L2_j_7,
	dbeta_L2,
	dalpha_L3_j_0, dalpha_L3_j_1, dalpha_L3_j_2, dalpha_L3_j_3, dalpha_L3_j_4,
	dbeta_L3,
	SIGN_dalpha_L1_j_0, SIGN_dalpha_L1_j_1, SIGN_dalpha_L1_j_2, SIGN_dalpha_L1_j_3, SIGN_dalpha_L1_j_4, SIGN_dalpha_L1_j_5, SIGN_dalpha_L1_j_6, SIGN_dalpha_L1_j_7, SIGN_dalpha_L1_j_8, SIGN_dalpha_L1_j_9, SIGN_dalpha_L1_j_10, SIGN_dalpha_L1_j_11, SIGN_dalpha_L1_j_12, SIGN_dalpha_L1_j_13, SIGN_dalpha_L1_j_14, SIGN_dalpha_L1_j_15, SIGN_dalpha_L1_j_16, SIGN_dalpha_L1_j_17, SIGN_dalpha_L1_j_18, SIGN_dalpha_L1_j_19, SIGN_dalpha_L1_j_20, SIGN_dalpha_L1_j_21, SIGN_dalpha_L1_j_22, SIGN_dalpha_L1_j_23, SIGN_dalpha_L1_j_24,
	SIGN_dbeta_L1,
	SIGN_dalpha_L2_j_0, SIGN_dalpha_L2_j_1, SIGN_dalpha_L2_j_2, SIGN_dalpha_L2_j_3, SIGN_dalpha_L2_j_4, SIGN_dalpha_L2_j_5, SIGN_dalpha_L2_j_6, SIGN_dalpha_L2_j_7,
	SIGN_dbeta_L2,
	SIGN_dalpha_L3_j_0, SIGN_dalpha_L3_j_1, SIGN_dalpha_L3_j_2, SIGN_dalpha_L3_j_3, SIGN_dalpha_L3_j_4,
	SIGN_dbeta_L3,
	rc,
	CLK, INIT
);

input wire [5 - 1:0] dalpha_L1_j_0_netPar0, dalpha_L1_j_1_netPar0, dalpha_L1_j_2_netPar0, dalpha_L1_j_3_netPar0, dalpha_L1_j_4_netPar0, dalpha_L1_j_5_netPar0, dalpha_L1_j_6_netPar0, dalpha_L1_j_7_netPar0, dalpha_L1_j_8_netPar0, dalpha_L1_j_9_netPar0, dalpha_L1_j_10_netPar0, dalpha_L1_j_11_netPar0, dalpha_L1_j_12_netPar0, dalpha_L1_j_13_netPar0, dalpha_L1_j_14_netPar0, dalpha_L1_j_15_netPar0, dalpha_L1_j_16_netPar0, dalpha_L1_j_17_netPar0, dalpha_L1_j_18_netPar0, dalpha_L1_j_19_netPar0, dalpha_L1_j_20_netPar0, dalpha_L1_j_21_netPar0, dalpha_L1_j_22_netPar0, dalpha_L1_j_23_netPar0, dalpha_L1_j_24_netPar0;
input wire [25 - 1:0] dbeta_L1_netPar0;
input wire [25 - 1:0] dalpha_L2_j_0_netPar0, dalpha_L2_j_1_netPar0, dalpha_L2_j_2_netPar0, dalpha_L2_j_3_netPar0, dalpha_L2_j_4_netPar0, dalpha_L2_j_5_netPar0, dalpha_L2_j_6_netPar0, dalpha_L2_j_7_netPar0;
input wire [8 - 1:0] dbeta_L2_netPar0;
input wire [8 - 1:0] dalpha_L3_j_0_netPar0, dalpha_L3_j_1_netPar0, dalpha_L3_j_2_netPar0, dalpha_L3_j_3_netPar0, dalpha_L3_j_4_netPar0;
input wire [5 - 1:0] dbeta_L3_netPar0;
input wire [5 - 1:0] SIGN_dalpha_L1_j_0_netPar0, SIGN_dalpha_L1_j_1_netPar0, SIGN_dalpha_L1_j_2_netPar0, SIGN_dalpha_L1_j_3_netPar0, SIGN_dalpha_L1_j_4_netPar0, SIGN_dalpha_L1_j_5_netPar0, SIGN_dalpha_L1_j_6_netPar0, SIGN_dalpha_L1_j_7_netPar0, SIGN_dalpha_L1_j_8_netPar0, SIGN_dalpha_L1_j_9_netPar0, SIGN_dalpha_L1_j_10_netPar0, SIGN_dalpha_L1_j_11_netPar0, SIGN_dalpha_L1_j_12_netPar0, SIGN_dalpha_L1_j_13_netPar0, SIGN_dalpha_L1_j_14_netPar0, SIGN_dalpha_L1_j_15_netPar0, SIGN_dalpha_L1_j_16_netPar0, SIGN_dalpha_L1_j_17_netPar0, SIGN_dalpha_L1_j_18_netPar0, SIGN_dalpha_L1_j_19_netPar0, SIGN_dalpha_L1_j_20_netPar0, SIGN_dalpha_L1_j_21_netPar0, SIGN_dalpha_L1_j_22_netPar0, SIGN_dalpha_L1_j_23_netPar0, SIGN_dalpha_L1_j_24_netPar0;
input wire [25 - 1:0] SIGN_dbeta_L1_netPar0;
input wire [25 - 1:0] SIGN_dalpha_L2_j_0_netPar0, SIGN_dalpha_L2_j_1_netPar0, SIGN_dalpha_L2_j_2_netPar0, SIGN_dalpha_L2_j_3_netPar0, SIGN_dalpha_L2_j_4_netPar0, SIGN_dalpha_L2_j_5_netPar0, SIGN_dalpha_L2_j_6_netPar0, SIGN_dalpha_L2_j_7_netPar0;
input wire [8 - 1:0] SIGN_dbeta_L2_netPar0;
input wire [8 - 1:0] SIGN_dalpha_L3_j_0_netPar0, SIGN_dalpha_L3_j_1_netPar0, SIGN_dalpha_L3_j_2_netPar0, SIGN_dalpha_L3_j_3_netPar0, SIGN_dalpha_L3_j_4_netPar0;
input wire [5 - 1:0] SIGN_dbeta_L3_netPar0;
input wire [5 - 1:0] dalpha_L1_j_0_netPar1, dalpha_L1_j_1_netPar1, dalpha_L1_j_2_netPar1, dalpha_L1_j_3_netPar1, dalpha_L1_j_4_netPar1, dalpha_L1_j_5_netPar1, dalpha_L1_j_6_netPar1, dalpha_L1_j_7_netPar1, dalpha_L1_j_8_netPar1, dalpha_L1_j_9_netPar1, dalpha_L1_j_10_netPar1, dalpha_L1_j_11_netPar1, dalpha_L1_j_12_netPar1, dalpha_L1_j_13_netPar1, dalpha_L1_j_14_netPar1, dalpha_L1_j_15_netPar1, dalpha_L1_j_16_netPar1, dalpha_L1_j_17_netPar1, dalpha_L1_j_18_netPar1, dalpha_L1_j_19_netPar1, dalpha_L1_j_20_netPar1, dalpha_L1_j_21_netPar1, dalpha_L1_j_22_netPar1, dalpha_L1_j_23_netPar1, dalpha_L1_j_24_netPar1;
input wire [25 - 1:0] dbeta_L1_netPar1;
input wire [25 - 1:0] dalpha_L2_j_0_netPar1, dalpha_L2_j_1_netPar1, dalpha_L2_j_2_netPar1, dalpha_L2_j_3_netPar1, dalpha_L2_j_4_netPar1, dalpha_L2_j_5_netPar1, dalpha_L2_j_6_netPar1, dalpha_L2_j_7_netPar1;
input wire [8 - 1:0] dbeta_L2_netPar1;
input wire [8 - 1:0] dalpha_L3_j_0_netPar1, dalpha_L3_j_1_netPar1, dalpha_L3_j_2_netPar1, dalpha_L3_j_3_netPar1, dalpha_L3_j_4_netPar1;
input wire [5 - 1:0] dbeta_L3_netPar1;
input wire [5 - 1:0] SIGN_dalpha_L1_j_0_netPar1, SIGN_dalpha_L1_j_1_netPar1, SIGN_dalpha_L1_j_2_netPar1, SIGN_dalpha_L1_j_3_netPar1, SIGN_dalpha_L1_j_4_netPar1, SIGN_dalpha_L1_j_5_netPar1, SIGN_dalpha_L1_j_6_netPar1, SIGN_dalpha_L1_j_7_netPar1, SIGN_dalpha_L1_j_8_netPar1, SIGN_dalpha_L1_j_9_netPar1, SIGN_dalpha_L1_j_10_netPar1, SIGN_dalpha_L1_j_11_netPar1, SIGN_dalpha_L1_j_12_netPar1, SIGN_dalpha_L1_j_13_netPar1, SIGN_dalpha_L1_j_14_netPar1, SIGN_dalpha_L1_j_15_netPar1, SIGN_dalpha_L1_j_16_netPar1, SIGN_dalpha_L1_j_17_netPar1, SIGN_dalpha_L1_j_18_netPar1, SIGN_dalpha_L1_j_19_netPar1, SIGN_dalpha_L1_j_20_netPar1, SIGN_dalpha_L1_j_21_netPar1, SIGN_dalpha_L1_j_22_netPar1, SIGN_dalpha_L1_j_23_netPar1, SIGN_dalpha_L1_j_24_netPar1;
input wire [25 - 1:0] SIGN_dbeta_L1_netPar1;
input wire [25 - 1:0] SIGN_dalpha_L2_j_0_netPar1, SIGN_dalpha_L2_j_1_netPar1, SIGN_dalpha_L2_j_2_netPar1, SIGN_dalpha_L2_j_3_netPar1, SIGN_dalpha_L2_j_4_netPar1, SIGN_dalpha_L2_j_5_netPar1, SIGN_dalpha_L2_j_6_netPar1, SIGN_dalpha_L2_j_7_netPar1;
input wire [8 - 1:0] SIGN_dbeta_L2_netPar1;
input wire [8 - 1:0] SIGN_dalpha_L3_j_0_netPar1, SIGN_dalpha_L3_j_1_netPar1, SIGN_dalpha_L3_j_2_netPar1, SIGN_dalpha_L3_j_3_netPar1, SIGN_dalpha_L3_j_4_netPar1;
input wire [5 - 1:0] SIGN_dbeta_L3_netPar1;
input wire [5 - 1:0] dalpha_L1_j_0_netPar2, dalpha_L1_j_1_netPar2, dalpha_L1_j_2_netPar2, dalpha_L1_j_3_netPar2, dalpha_L1_j_4_netPar2, dalpha_L1_j_5_netPar2, dalpha_L1_j_6_netPar2, dalpha_L1_j_7_netPar2, dalpha_L1_j_8_netPar2, dalpha_L1_j_9_netPar2, dalpha_L1_j_10_netPar2, dalpha_L1_j_11_netPar2, dalpha_L1_j_12_netPar2, dalpha_L1_j_13_netPar2, dalpha_L1_j_14_netPar2, dalpha_L1_j_15_netPar2, dalpha_L1_j_16_netPar2, dalpha_L1_j_17_netPar2, dalpha_L1_j_18_netPar2, dalpha_L1_j_19_netPar2, dalpha_L1_j_20_netPar2, dalpha_L1_j_21_netPar2, dalpha_L1_j_22_netPar2, dalpha_L1_j_23_netPar2, dalpha_L1_j_24_netPar2;
input wire [25 - 1:0] dbeta_L1_netPar2;
input wire [25 - 1:0] dalpha_L2_j_0_netPar2, dalpha_L2_j_1_netPar2, dalpha_L2_j_2_netPar2, dalpha_L2_j_3_netPar2, dalpha_L2_j_4_netPar2, dalpha_L2_j_5_netPar2, dalpha_L2_j_6_netPar2, dalpha_L2_j_7_netPar2;
input wire [8 - 1:0] dbeta_L2_netPar2;
input wire [8 - 1:0] dalpha_L3_j_0_netPar2, dalpha_L3_j_1_netPar2, dalpha_L3_j_2_netPar2, dalpha_L3_j_3_netPar2, dalpha_L3_j_4_netPar2;
input wire [5 - 1:0] dbeta_L3_netPar2;
input wire [5 - 1:0] SIGN_dalpha_L1_j_0_netPar2, SIGN_dalpha_L1_j_1_netPar2, SIGN_dalpha_L1_j_2_netPar2, SIGN_dalpha_L1_j_3_netPar2, SIGN_dalpha_L1_j_4_netPar2, SIGN_dalpha_L1_j_5_netPar2, SIGN_dalpha_L1_j_6_netPar2, SIGN_dalpha_L1_j_7_netPar2, SIGN_dalpha_L1_j_8_netPar2, SIGN_dalpha_L1_j_9_netPar2, SIGN_dalpha_L1_j_10_netPar2, SIGN_dalpha_L1_j_11_netPar2, SIGN_dalpha_L1_j_12_netPar2, SIGN_dalpha_L1_j_13_netPar2, SIGN_dalpha_L1_j_14_netPar2, SIGN_dalpha_L1_j_15_netPar2, SIGN_dalpha_L1_j_16_netPar2, SIGN_dalpha_L1_j_17_netPar2, SIGN_dalpha_L1_j_18_netPar2, SIGN_dalpha_L1_j_19_netPar2, SIGN_dalpha_L1_j_20_netPar2, SIGN_dalpha_L1_j_21_netPar2, SIGN_dalpha_L1_j_22_netPar2, SIGN_dalpha_L1_j_23_netPar2, SIGN_dalpha_L1_j_24_netPar2;
input wire [25 - 1:0] SIGN_dbeta_L1_netPar2;
input wire [25 - 1:0] SIGN_dalpha_L2_j_0_netPar2, SIGN_dalpha_L2_j_1_netPar2, SIGN_dalpha_L2_j_2_netPar2, SIGN_dalpha_L2_j_3_netPar2, SIGN_dalpha_L2_j_4_netPar2, SIGN_dalpha_L2_j_5_netPar2, SIGN_dalpha_L2_j_6_netPar2, SIGN_dalpha_L2_j_7_netPar2;
input wire [8 - 1:0] SIGN_dbeta_L2_netPar2;
input wire [8 - 1:0] SIGN_dalpha_L3_j_0_netPar2, SIGN_dalpha_L3_j_1_netPar2, SIGN_dalpha_L3_j_2_netPar2, SIGN_dalpha_L3_j_3_netPar2, SIGN_dalpha_L3_j_4_netPar2;
input wire [5 - 1:0] SIGN_dbeta_L3_netPar2;

input wire [408-1:0] rc;

input wire CLK, INIT;

output wire [5 - 1:0] dalpha_L1_j_0, dalpha_L1_j_1, dalpha_L1_j_2, dalpha_L1_j_3, dalpha_L1_j_4, dalpha_L1_j_5, dalpha_L1_j_6, dalpha_L1_j_7, dalpha_L1_j_8, dalpha_L1_j_9, dalpha_L1_j_10, dalpha_L1_j_11, dalpha_L1_j_12, dalpha_L1_j_13, dalpha_L1_j_14, dalpha_L1_j_15, dalpha_L1_j_16, dalpha_L1_j_17, dalpha_L1_j_18, dalpha_L1_j_19, dalpha_L1_j_20, dalpha_L1_j_21, dalpha_L1_j_22, dalpha_L1_j_23, dalpha_L1_j_24;
output wire [25 - 1:0] dbeta_L1;
output wire [25 - 1:0] dalpha_L2_j_0, dalpha_L2_j_1, dalpha_L2_j_2, dalpha_L2_j_3, dalpha_L2_j_4, dalpha_L2_j_5, dalpha_L2_j_6, dalpha_L2_j_7;
output wire [8 - 1:0] dbeta_L2;
output wire [8 - 1:0] dalpha_L3_j_0, dalpha_L3_j_1, dalpha_L3_j_2, dalpha_L3_j_3, dalpha_L3_j_4;
output wire [5 - 1:0] dbeta_L3;
output wire [5 - 1:0] SIGN_dalpha_L1_j_0, SIGN_dalpha_L1_j_1, SIGN_dalpha_L1_j_2, SIGN_dalpha_L1_j_3, SIGN_dalpha_L1_j_4, SIGN_dalpha_L1_j_5, SIGN_dalpha_L1_j_6, SIGN_dalpha_L1_j_7, SIGN_dalpha_L1_j_8, SIGN_dalpha_L1_j_9, SIGN_dalpha_L1_j_10, SIGN_dalpha_L1_j_11, SIGN_dalpha_L1_j_12, SIGN_dalpha_L1_j_13, SIGN_dalpha_L1_j_14, SIGN_dalpha_L1_j_15, SIGN_dalpha_L1_j_16, SIGN_dalpha_L1_j_17, SIGN_dalpha_L1_j_18, SIGN_dalpha_L1_j_19, SIGN_dalpha_L1_j_20, SIGN_dalpha_L1_j_21, SIGN_dalpha_L1_j_22, SIGN_dalpha_L1_j_23, SIGN_dalpha_L1_j_24;
output wire [25 - 1:0] SIGN_dbeta_L1;
output wire [25 - 1:0] SIGN_dalpha_L2_j_0, SIGN_dalpha_L2_j_1, SIGN_dalpha_L2_j_2, SIGN_dalpha_L2_j_3, SIGN_dalpha_L2_j_4, SIGN_dalpha_L2_j_5, SIGN_dalpha_L2_j_6, SIGN_dalpha_L2_j_7;
output wire [8 - 1:0] SIGN_dbeta_L2;
output wire [8 - 1:0] SIGN_dalpha_L3_j_0, SIGN_dalpha_L3_j_1, SIGN_dalpha_L3_j_2, SIGN_dalpha_L3_j_3, SIGN_dalpha_L3_j_4;
output wire [5 - 1:0] SIGN_dbeta_L3;

SS_ADDSUB ADDSUB_dalpha_L1_0_0(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_0_netPar0[0], dalpha_L1_j_0_netPar1[0], dalpha_L1_j_0_netPar2[0] }), .SIGN({ SIGN_dalpha_L1_j_0_netPar0[0], SIGN_dalpha_L1_j_0_netPar1[0], SIGN_dalpha_L1_j_0_netPar2[0]}), .R_condition(rc[0]), .OUT(dalpha_L1_j_0[0]), .SIGN_out(SIGN_dalpha_L1_j_0[0]));
SS_ADDSUB ADDSUB_dalpha_L1_0_1(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_1_netPar0[0], dalpha_L1_j_1_netPar1[0], dalpha_L1_j_1_netPar2[0] }), .SIGN({ SIGN_dalpha_L1_j_1_netPar0[0], SIGN_dalpha_L1_j_1_netPar1[0], SIGN_dalpha_L1_j_1_netPar2[0]}), .R_condition(rc[1]), .OUT(dalpha_L1_j_1[0]), .SIGN_out(SIGN_dalpha_L1_j_1[0]));
SS_ADDSUB ADDSUB_dalpha_L1_0_2(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_2_netPar0[0], dalpha_L1_j_2_netPar1[0], dalpha_L1_j_2_netPar2[0] }), .SIGN({ SIGN_dalpha_L1_j_2_netPar0[0], SIGN_dalpha_L1_j_2_netPar1[0], SIGN_dalpha_L1_j_2_netPar2[0]}), .R_condition(rc[2]), .OUT(dalpha_L1_j_2[0]), .SIGN_out(SIGN_dalpha_L1_j_2[0]));
SS_ADDSUB ADDSUB_dalpha_L1_0_3(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_3_netPar0[0], dalpha_L1_j_3_netPar1[0], dalpha_L1_j_3_netPar2[0] }), .SIGN({ SIGN_dalpha_L1_j_3_netPar0[0], SIGN_dalpha_L1_j_3_netPar1[0], SIGN_dalpha_L1_j_3_netPar2[0]}), .R_condition(rc[3]), .OUT(dalpha_L1_j_3[0]), .SIGN_out(SIGN_dalpha_L1_j_3[0]));
SS_ADDSUB ADDSUB_dalpha_L1_0_4(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_4_netPar0[0], dalpha_L1_j_4_netPar1[0], dalpha_L1_j_4_netPar2[0] }), .SIGN({ SIGN_dalpha_L1_j_4_netPar0[0], SIGN_dalpha_L1_j_4_netPar1[0], SIGN_dalpha_L1_j_4_netPar2[0]}), .R_condition(rc[4]), .OUT(dalpha_L1_j_4[0]), .SIGN_out(SIGN_dalpha_L1_j_4[0]));
SS_ADDSUB ADDSUB_dalpha_L1_0_5(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_5_netPar0[0], dalpha_L1_j_5_netPar1[0], dalpha_L1_j_5_netPar2[0] }), .SIGN({ SIGN_dalpha_L1_j_5_netPar0[0], SIGN_dalpha_L1_j_5_netPar1[0], SIGN_dalpha_L1_j_5_netPar2[0]}), .R_condition(rc[5]), .OUT(dalpha_L1_j_5[0]), .SIGN_out(SIGN_dalpha_L1_j_5[0]));
SS_ADDSUB ADDSUB_dalpha_L1_0_6(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_6_netPar0[0], dalpha_L1_j_6_netPar1[0], dalpha_L1_j_6_netPar2[0] }), .SIGN({ SIGN_dalpha_L1_j_6_netPar0[0], SIGN_dalpha_L1_j_6_netPar1[0], SIGN_dalpha_L1_j_6_netPar2[0]}), .R_condition(rc[6]), .OUT(dalpha_L1_j_6[0]), .SIGN_out(SIGN_dalpha_L1_j_6[0]));
SS_ADDSUB ADDSUB_dalpha_L1_0_7(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_7_netPar0[0], dalpha_L1_j_7_netPar1[0], dalpha_L1_j_7_netPar2[0] }), .SIGN({ SIGN_dalpha_L1_j_7_netPar0[0], SIGN_dalpha_L1_j_7_netPar1[0], SIGN_dalpha_L1_j_7_netPar2[0]}), .R_condition(rc[7]), .OUT(dalpha_L1_j_7[0]), .SIGN_out(SIGN_dalpha_L1_j_7[0]));
SS_ADDSUB ADDSUB_dalpha_L1_0_8(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_8_netPar0[0], dalpha_L1_j_8_netPar1[0], dalpha_L1_j_8_netPar2[0] }), .SIGN({ SIGN_dalpha_L1_j_8_netPar0[0], SIGN_dalpha_L1_j_8_netPar1[0], SIGN_dalpha_L1_j_8_netPar2[0]}), .R_condition(rc[8]), .OUT(dalpha_L1_j_8[0]), .SIGN_out(SIGN_dalpha_L1_j_8[0]));
SS_ADDSUB ADDSUB_dalpha_L1_0_9(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_9_netPar0[0], dalpha_L1_j_9_netPar1[0], dalpha_L1_j_9_netPar2[0] }), .SIGN({ SIGN_dalpha_L1_j_9_netPar0[0], SIGN_dalpha_L1_j_9_netPar1[0], SIGN_dalpha_L1_j_9_netPar2[0]}), .R_condition(rc[9]), .OUT(dalpha_L1_j_9[0]), .SIGN_out(SIGN_dalpha_L1_j_9[0]));
SS_ADDSUB ADDSUB_dalpha_L1_0_10(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_10_netPar0[0], dalpha_L1_j_10_netPar1[0], dalpha_L1_j_10_netPar2[0] }), .SIGN({ SIGN_dalpha_L1_j_10_netPar0[0], SIGN_dalpha_L1_j_10_netPar1[0], SIGN_dalpha_L1_j_10_netPar2[0]}), .R_condition(rc[10]), .OUT(dalpha_L1_j_10[0]), .SIGN_out(SIGN_dalpha_L1_j_10[0]));
SS_ADDSUB ADDSUB_dalpha_L1_0_11(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_11_netPar0[0], dalpha_L1_j_11_netPar1[0], dalpha_L1_j_11_netPar2[0] }), .SIGN({ SIGN_dalpha_L1_j_11_netPar0[0], SIGN_dalpha_L1_j_11_netPar1[0], SIGN_dalpha_L1_j_11_netPar2[0]}), .R_condition(rc[11]), .OUT(dalpha_L1_j_11[0]), .SIGN_out(SIGN_dalpha_L1_j_11[0]));
SS_ADDSUB ADDSUB_dalpha_L1_0_12(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_12_netPar0[0], dalpha_L1_j_12_netPar1[0], dalpha_L1_j_12_netPar2[0] }), .SIGN({ SIGN_dalpha_L1_j_12_netPar0[0], SIGN_dalpha_L1_j_12_netPar1[0], SIGN_dalpha_L1_j_12_netPar2[0]}), .R_condition(rc[12]), .OUT(dalpha_L1_j_12[0]), .SIGN_out(SIGN_dalpha_L1_j_12[0]));
SS_ADDSUB ADDSUB_dalpha_L1_0_13(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_13_netPar0[0], dalpha_L1_j_13_netPar1[0], dalpha_L1_j_13_netPar2[0] }), .SIGN({ SIGN_dalpha_L1_j_13_netPar0[0], SIGN_dalpha_L1_j_13_netPar1[0], SIGN_dalpha_L1_j_13_netPar2[0]}), .R_condition(rc[13]), .OUT(dalpha_L1_j_13[0]), .SIGN_out(SIGN_dalpha_L1_j_13[0]));
SS_ADDSUB ADDSUB_dalpha_L1_0_14(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_14_netPar0[0], dalpha_L1_j_14_netPar1[0], dalpha_L1_j_14_netPar2[0] }), .SIGN({ SIGN_dalpha_L1_j_14_netPar0[0], SIGN_dalpha_L1_j_14_netPar1[0], SIGN_dalpha_L1_j_14_netPar2[0]}), .R_condition(rc[14]), .OUT(dalpha_L1_j_14[0]), .SIGN_out(SIGN_dalpha_L1_j_14[0]));
SS_ADDSUB ADDSUB_dalpha_L1_0_15(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_15_netPar0[0], dalpha_L1_j_15_netPar1[0], dalpha_L1_j_15_netPar2[0] }), .SIGN({ SIGN_dalpha_L1_j_15_netPar0[0], SIGN_dalpha_L1_j_15_netPar1[0], SIGN_dalpha_L1_j_15_netPar2[0]}), .R_condition(rc[15]), .OUT(dalpha_L1_j_15[0]), .SIGN_out(SIGN_dalpha_L1_j_15[0]));
SS_ADDSUB ADDSUB_dalpha_L1_0_16(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_16_netPar0[0], dalpha_L1_j_16_netPar1[0], dalpha_L1_j_16_netPar2[0] }), .SIGN({ SIGN_dalpha_L1_j_16_netPar0[0], SIGN_dalpha_L1_j_16_netPar1[0], SIGN_dalpha_L1_j_16_netPar2[0]}), .R_condition(rc[16]), .OUT(dalpha_L1_j_16[0]), .SIGN_out(SIGN_dalpha_L1_j_16[0]));
SS_ADDSUB ADDSUB_dalpha_L1_0_17(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_17_netPar0[0], dalpha_L1_j_17_netPar1[0], dalpha_L1_j_17_netPar2[0] }), .SIGN({ SIGN_dalpha_L1_j_17_netPar0[0], SIGN_dalpha_L1_j_17_netPar1[0], SIGN_dalpha_L1_j_17_netPar2[0]}), .R_condition(rc[17]), .OUT(dalpha_L1_j_17[0]), .SIGN_out(SIGN_dalpha_L1_j_17[0]));
SS_ADDSUB ADDSUB_dalpha_L1_0_18(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_18_netPar0[0], dalpha_L1_j_18_netPar1[0], dalpha_L1_j_18_netPar2[0] }), .SIGN({ SIGN_dalpha_L1_j_18_netPar0[0], SIGN_dalpha_L1_j_18_netPar1[0], SIGN_dalpha_L1_j_18_netPar2[0]}), .R_condition(rc[18]), .OUT(dalpha_L1_j_18[0]), .SIGN_out(SIGN_dalpha_L1_j_18[0]));
SS_ADDSUB ADDSUB_dalpha_L1_0_19(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_19_netPar0[0], dalpha_L1_j_19_netPar1[0], dalpha_L1_j_19_netPar2[0] }), .SIGN({ SIGN_dalpha_L1_j_19_netPar0[0], SIGN_dalpha_L1_j_19_netPar1[0], SIGN_dalpha_L1_j_19_netPar2[0]}), .R_condition(rc[19]), .OUT(dalpha_L1_j_19[0]), .SIGN_out(SIGN_dalpha_L1_j_19[0]));
SS_ADDSUB ADDSUB_dalpha_L1_0_20(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_20_netPar0[0], dalpha_L1_j_20_netPar1[0], dalpha_L1_j_20_netPar2[0] }), .SIGN({ SIGN_dalpha_L1_j_20_netPar0[0], SIGN_dalpha_L1_j_20_netPar1[0], SIGN_dalpha_L1_j_20_netPar2[0]}), .R_condition(rc[20]), .OUT(dalpha_L1_j_20[0]), .SIGN_out(SIGN_dalpha_L1_j_20[0]));
SS_ADDSUB ADDSUB_dalpha_L1_0_21(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_21_netPar0[0], dalpha_L1_j_21_netPar1[0], dalpha_L1_j_21_netPar2[0] }), .SIGN({ SIGN_dalpha_L1_j_21_netPar0[0], SIGN_dalpha_L1_j_21_netPar1[0], SIGN_dalpha_L1_j_21_netPar2[0]}), .R_condition(rc[21]), .OUT(dalpha_L1_j_21[0]), .SIGN_out(SIGN_dalpha_L1_j_21[0]));
SS_ADDSUB ADDSUB_dalpha_L1_0_22(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_22_netPar0[0], dalpha_L1_j_22_netPar1[0], dalpha_L1_j_22_netPar2[0] }), .SIGN({ SIGN_dalpha_L1_j_22_netPar0[0], SIGN_dalpha_L1_j_22_netPar1[0], SIGN_dalpha_L1_j_22_netPar2[0]}), .R_condition(rc[22]), .OUT(dalpha_L1_j_22[0]), .SIGN_out(SIGN_dalpha_L1_j_22[0]));
SS_ADDSUB ADDSUB_dalpha_L1_0_23(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_23_netPar0[0], dalpha_L1_j_23_netPar1[0], dalpha_L1_j_23_netPar2[0] }), .SIGN({ SIGN_dalpha_L1_j_23_netPar0[0], SIGN_dalpha_L1_j_23_netPar1[0], SIGN_dalpha_L1_j_23_netPar2[0]}), .R_condition(rc[23]), .OUT(dalpha_L1_j_23[0]), .SIGN_out(SIGN_dalpha_L1_j_23[0]));
SS_ADDSUB ADDSUB_dalpha_L1_0_24(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_24_netPar0[0], dalpha_L1_j_24_netPar1[0], dalpha_L1_j_24_netPar2[0] }), .SIGN({ SIGN_dalpha_L1_j_24_netPar0[0], SIGN_dalpha_L1_j_24_netPar1[0], SIGN_dalpha_L1_j_24_netPar2[0]}), .R_condition(rc[24]), .OUT(dalpha_L1_j_24[0]), .SIGN_out(SIGN_dalpha_L1_j_24[0]));
SS_ADDSUB ADDSUB_dalpha_L1_1_0(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_0_netPar0[1], dalpha_L1_j_0_netPar1[1], dalpha_L1_j_0_netPar2[1] }), .SIGN({ SIGN_dalpha_L1_j_0_netPar0[1], SIGN_dalpha_L1_j_0_netPar1[1], SIGN_dalpha_L1_j_0_netPar2[1]}), .R_condition(rc[25]), .OUT(dalpha_L1_j_0[1]), .SIGN_out(SIGN_dalpha_L1_j_0[1]));
SS_ADDSUB ADDSUB_dalpha_L1_1_1(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_1_netPar0[1], dalpha_L1_j_1_netPar1[1], dalpha_L1_j_1_netPar2[1] }), .SIGN({ SIGN_dalpha_L1_j_1_netPar0[1], SIGN_dalpha_L1_j_1_netPar1[1], SIGN_dalpha_L1_j_1_netPar2[1]}), .R_condition(rc[26]), .OUT(dalpha_L1_j_1[1]), .SIGN_out(SIGN_dalpha_L1_j_1[1]));
SS_ADDSUB ADDSUB_dalpha_L1_1_2(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_2_netPar0[1], dalpha_L1_j_2_netPar1[1], dalpha_L1_j_2_netPar2[1] }), .SIGN({ SIGN_dalpha_L1_j_2_netPar0[1], SIGN_dalpha_L1_j_2_netPar1[1], SIGN_dalpha_L1_j_2_netPar2[1]}), .R_condition(rc[27]), .OUT(dalpha_L1_j_2[1]), .SIGN_out(SIGN_dalpha_L1_j_2[1]));
SS_ADDSUB ADDSUB_dalpha_L1_1_3(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_3_netPar0[1], dalpha_L1_j_3_netPar1[1], dalpha_L1_j_3_netPar2[1] }), .SIGN({ SIGN_dalpha_L1_j_3_netPar0[1], SIGN_dalpha_L1_j_3_netPar1[1], SIGN_dalpha_L1_j_3_netPar2[1]}), .R_condition(rc[28]), .OUT(dalpha_L1_j_3[1]), .SIGN_out(SIGN_dalpha_L1_j_3[1]));
SS_ADDSUB ADDSUB_dalpha_L1_1_4(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_4_netPar0[1], dalpha_L1_j_4_netPar1[1], dalpha_L1_j_4_netPar2[1] }), .SIGN({ SIGN_dalpha_L1_j_4_netPar0[1], SIGN_dalpha_L1_j_4_netPar1[1], SIGN_dalpha_L1_j_4_netPar2[1]}), .R_condition(rc[29]), .OUT(dalpha_L1_j_4[1]), .SIGN_out(SIGN_dalpha_L1_j_4[1]));
SS_ADDSUB ADDSUB_dalpha_L1_1_5(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_5_netPar0[1], dalpha_L1_j_5_netPar1[1], dalpha_L1_j_5_netPar2[1] }), .SIGN({ SIGN_dalpha_L1_j_5_netPar0[1], SIGN_dalpha_L1_j_5_netPar1[1], SIGN_dalpha_L1_j_5_netPar2[1]}), .R_condition(rc[30]), .OUT(dalpha_L1_j_5[1]), .SIGN_out(SIGN_dalpha_L1_j_5[1]));
SS_ADDSUB ADDSUB_dalpha_L1_1_6(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_6_netPar0[1], dalpha_L1_j_6_netPar1[1], dalpha_L1_j_6_netPar2[1] }), .SIGN({ SIGN_dalpha_L1_j_6_netPar0[1], SIGN_dalpha_L1_j_6_netPar1[1], SIGN_dalpha_L1_j_6_netPar2[1]}), .R_condition(rc[31]), .OUT(dalpha_L1_j_6[1]), .SIGN_out(SIGN_dalpha_L1_j_6[1]));
SS_ADDSUB ADDSUB_dalpha_L1_1_7(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_7_netPar0[1], dalpha_L1_j_7_netPar1[1], dalpha_L1_j_7_netPar2[1] }), .SIGN({ SIGN_dalpha_L1_j_7_netPar0[1], SIGN_dalpha_L1_j_7_netPar1[1], SIGN_dalpha_L1_j_7_netPar2[1]}), .R_condition(rc[32]), .OUT(dalpha_L1_j_7[1]), .SIGN_out(SIGN_dalpha_L1_j_7[1]));
SS_ADDSUB ADDSUB_dalpha_L1_1_8(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_8_netPar0[1], dalpha_L1_j_8_netPar1[1], dalpha_L1_j_8_netPar2[1] }), .SIGN({ SIGN_dalpha_L1_j_8_netPar0[1], SIGN_dalpha_L1_j_8_netPar1[1], SIGN_dalpha_L1_j_8_netPar2[1]}), .R_condition(rc[33]), .OUT(dalpha_L1_j_8[1]), .SIGN_out(SIGN_dalpha_L1_j_8[1]));
SS_ADDSUB ADDSUB_dalpha_L1_1_9(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_9_netPar0[1], dalpha_L1_j_9_netPar1[1], dalpha_L1_j_9_netPar2[1] }), .SIGN({ SIGN_dalpha_L1_j_9_netPar0[1], SIGN_dalpha_L1_j_9_netPar1[1], SIGN_dalpha_L1_j_9_netPar2[1]}), .R_condition(rc[34]), .OUT(dalpha_L1_j_9[1]), .SIGN_out(SIGN_dalpha_L1_j_9[1]));
SS_ADDSUB ADDSUB_dalpha_L1_1_10(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_10_netPar0[1], dalpha_L1_j_10_netPar1[1], dalpha_L1_j_10_netPar2[1] }), .SIGN({ SIGN_dalpha_L1_j_10_netPar0[1], SIGN_dalpha_L1_j_10_netPar1[1], SIGN_dalpha_L1_j_10_netPar2[1]}), .R_condition(rc[35]), .OUT(dalpha_L1_j_10[1]), .SIGN_out(SIGN_dalpha_L1_j_10[1]));
SS_ADDSUB ADDSUB_dalpha_L1_1_11(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_11_netPar0[1], dalpha_L1_j_11_netPar1[1], dalpha_L1_j_11_netPar2[1] }), .SIGN({ SIGN_dalpha_L1_j_11_netPar0[1], SIGN_dalpha_L1_j_11_netPar1[1], SIGN_dalpha_L1_j_11_netPar2[1]}), .R_condition(rc[36]), .OUT(dalpha_L1_j_11[1]), .SIGN_out(SIGN_dalpha_L1_j_11[1]));
SS_ADDSUB ADDSUB_dalpha_L1_1_12(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_12_netPar0[1], dalpha_L1_j_12_netPar1[1], dalpha_L1_j_12_netPar2[1] }), .SIGN({ SIGN_dalpha_L1_j_12_netPar0[1], SIGN_dalpha_L1_j_12_netPar1[1], SIGN_dalpha_L1_j_12_netPar2[1]}), .R_condition(rc[37]), .OUT(dalpha_L1_j_12[1]), .SIGN_out(SIGN_dalpha_L1_j_12[1]));
SS_ADDSUB ADDSUB_dalpha_L1_1_13(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_13_netPar0[1], dalpha_L1_j_13_netPar1[1], dalpha_L1_j_13_netPar2[1] }), .SIGN({ SIGN_dalpha_L1_j_13_netPar0[1], SIGN_dalpha_L1_j_13_netPar1[1], SIGN_dalpha_L1_j_13_netPar2[1]}), .R_condition(rc[38]), .OUT(dalpha_L1_j_13[1]), .SIGN_out(SIGN_dalpha_L1_j_13[1]));
SS_ADDSUB ADDSUB_dalpha_L1_1_14(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_14_netPar0[1], dalpha_L1_j_14_netPar1[1], dalpha_L1_j_14_netPar2[1] }), .SIGN({ SIGN_dalpha_L1_j_14_netPar0[1], SIGN_dalpha_L1_j_14_netPar1[1], SIGN_dalpha_L1_j_14_netPar2[1]}), .R_condition(rc[39]), .OUT(dalpha_L1_j_14[1]), .SIGN_out(SIGN_dalpha_L1_j_14[1]));
SS_ADDSUB ADDSUB_dalpha_L1_1_15(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_15_netPar0[1], dalpha_L1_j_15_netPar1[1], dalpha_L1_j_15_netPar2[1] }), .SIGN({ SIGN_dalpha_L1_j_15_netPar0[1], SIGN_dalpha_L1_j_15_netPar1[1], SIGN_dalpha_L1_j_15_netPar2[1]}), .R_condition(rc[40]), .OUT(dalpha_L1_j_15[1]), .SIGN_out(SIGN_dalpha_L1_j_15[1]));
SS_ADDSUB ADDSUB_dalpha_L1_1_16(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_16_netPar0[1], dalpha_L1_j_16_netPar1[1], dalpha_L1_j_16_netPar2[1] }), .SIGN({ SIGN_dalpha_L1_j_16_netPar0[1], SIGN_dalpha_L1_j_16_netPar1[1], SIGN_dalpha_L1_j_16_netPar2[1]}), .R_condition(rc[41]), .OUT(dalpha_L1_j_16[1]), .SIGN_out(SIGN_dalpha_L1_j_16[1]));
SS_ADDSUB ADDSUB_dalpha_L1_1_17(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_17_netPar0[1], dalpha_L1_j_17_netPar1[1], dalpha_L1_j_17_netPar2[1] }), .SIGN({ SIGN_dalpha_L1_j_17_netPar0[1], SIGN_dalpha_L1_j_17_netPar1[1], SIGN_dalpha_L1_j_17_netPar2[1]}), .R_condition(rc[42]), .OUT(dalpha_L1_j_17[1]), .SIGN_out(SIGN_dalpha_L1_j_17[1]));
SS_ADDSUB ADDSUB_dalpha_L1_1_18(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_18_netPar0[1], dalpha_L1_j_18_netPar1[1], dalpha_L1_j_18_netPar2[1] }), .SIGN({ SIGN_dalpha_L1_j_18_netPar0[1], SIGN_dalpha_L1_j_18_netPar1[1], SIGN_dalpha_L1_j_18_netPar2[1]}), .R_condition(rc[43]), .OUT(dalpha_L1_j_18[1]), .SIGN_out(SIGN_dalpha_L1_j_18[1]));
SS_ADDSUB ADDSUB_dalpha_L1_1_19(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_19_netPar0[1], dalpha_L1_j_19_netPar1[1], dalpha_L1_j_19_netPar2[1] }), .SIGN({ SIGN_dalpha_L1_j_19_netPar0[1], SIGN_dalpha_L1_j_19_netPar1[1], SIGN_dalpha_L1_j_19_netPar2[1]}), .R_condition(rc[44]), .OUT(dalpha_L1_j_19[1]), .SIGN_out(SIGN_dalpha_L1_j_19[1]));
SS_ADDSUB ADDSUB_dalpha_L1_1_20(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_20_netPar0[1], dalpha_L1_j_20_netPar1[1], dalpha_L1_j_20_netPar2[1] }), .SIGN({ SIGN_dalpha_L1_j_20_netPar0[1], SIGN_dalpha_L1_j_20_netPar1[1], SIGN_dalpha_L1_j_20_netPar2[1]}), .R_condition(rc[45]), .OUT(dalpha_L1_j_20[1]), .SIGN_out(SIGN_dalpha_L1_j_20[1]));
SS_ADDSUB ADDSUB_dalpha_L1_1_21(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_21_netPar0[1], dalpha_L1_j_21_netPar1[1], dalpha_L1_j_21_netPar2[1] }), .SIGN({ SIGN_dalpha_L1_j_21_netPar0[1], SIGN_dalpha_L1_j_21_netPar1[1], SIGN_dalpha_L1_j_21_netPar2[1]}), .R_condition(rc[46]), .OUT(dalpha_L1_j_21[1]), .SIGN_out(SIGN_dalpha_L1_j_21[1]));
SS_ADDSUB ADDSUB_dalpha_L1_1_22(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_22_netPar0[1], dalpha_L1_j_22_netPar1[1], dalpha_L1_j_22_netPar2[1] }), .SIGN({ SIGN_dalpha_L1_j_22_netPar0[1], SIGN_dalpha_L1_j_22_netPar1[1], SIGN_dalpha_L1_j_22_netPar2[1]}), .R_condition(rc[47]), .OUT(dalpha_L1_j_22[1]), .SIGN_out(SIGN_dalpha_L1_j_22[1]));
SS_ADDSUB ADDSUB_dalpha_L1_1_23(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_23_netPar0[1], dalpha_L1_j_23_netPar1[1], dalpha_L1_j_23_netPar2[1] }), .SIGN({ SIGN_dalpha_L1_j_23_netPar0[1], SIGN_dalpha_L1_j_23_netPar1[1], SIGN_dalpha_L1_j_23_netPar2[1]}), .R_condition(rc[48]), .OUT(dalpha_L1_j_23[1]), .SIGN_out(SIGN_dalpha_L1_j_23[1]));
SS_ADDSUB ADDSUB_dalpha_L1_1_24(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_24_netPar0[1], dalpha_L1_j_24_netPar1[1], dalpha_L1_j_24_netPar2[1] }), .SIGN({ SIGN_dalpha_L1_j_24_netPar0[1], SIGN_dalpha_L1_j_24_netPar1[1], SIGN_dalpha_L1_j_24_netPar2[1]}), .R_condition(rc[49]), .OUT(dalpha_L1_j_24[1]), .SIGN_out(SIGN_dalpha_L1_j_24[1]));
SS_ADDSUB ADDSUB_dalpha_L1_2_0(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_0_netPar0[2], dalpha_L1_j_0_netPar1[2], dalpha_L1_j_0_netPar2[2] }), .SIGN({ SIGN_dalpha_L1_j_0_netPar0[2], SIGN_dalpha_L1_j_0_netPar1[2], SIGN_dalpha_L1_j_0_netPar2[2]}), .R_condition(rc[50]), .OUT(dalpha_L1_j_0[2]), .SIGN_out(SIGN_dalpha_L1_j_0[2]));
SS_ADDSUB ADDSUB_dalpha_L1_2_1(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_1_netPar0[2], dalpha_L1_j_1_netPar1[2], dalpha_L1_j_1_netPar2[2] }), .SIGN({ SIGN_dalpha_L1_j_1_netPar0[2], SIGN_dalpha_L1_j_1_netPar1[2], SIGN_dalpha_L1_j_1_netPar2[2]}), .R_condition(rc[51]), .OUT(dalpha_L1_j_1[2]), .SIGN_out(SIGN_dalpha_L1_j_1[2]));
SS_ADDSUB ADDSUB_dalpha_L1_2_2(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_2_netPar0[2], dalpha_L1_j_2_netPar1[2], dalpha_L1_j_2_netPar2[2] }), .SIGN({ SIGN_dalpha_L1_j_2_netPar0[2], SIGN_dalpha_L1_j_2_netPar1[2], SIGN_dalpha_L1_j_2_netPar2[2]}), .R_condition(rc[52]), .OUT(dalpha_L1_j_2[2]), .SIGN_out(SIGN_dalpha_L1_j_2[2]));
SS_ADDSUB ADDSUB_dalpha_L1_2_3(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_3_netPar0[2], dalpha_L1_j_3_netPar1[2], dalpha_L1_j_3_netPar2[2] }), .SIGN({ SIGN_dalpha_L1_j_3_netPar0[2], SIGN_dalpha_L1_j_3_netPar1[2], SIGN_dalpha_L1_j_3_netPar2[2]}), .R_condition(rc[53]), .OUT(dalpha_L1_j_3[2]), .SIGN_out(SIGN_dalpha_L1_j_3[2]));
SS_ADDSUB ADDSUB_dalpha_L1_2_4(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_4_netPar0[2], dalpha_L1_j_4_netPar1[2], dalpha_L1_j_4_netPar2[2] }), .SIGN({ SIGN_dalpha_L1_j_4_netPar0[2], SIGN_dalpha_L1_j_4_netPar1[2], SIGN_dalpha_L1_j_4_netPar2[2]}), .R_condition(rc[54]), .OUT(dalpha_L1_j_4[2]), .SIGN_out(SIGN_dalpha_L1_j_4[2]));
SS_ADDSUB ADDSUB_dalpha_L1_2_5(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_5_netPar0[2], dalpha_L1_j_5_netPar1[2], dalpha_L1_j_5_netPar2[2] }), .SIGN({ SIGN_dalpha_L1_j_5_netPar0[2], SIGN_dalpha_L1_j_5_netPar1[2], SIGN_dalpha_L1_j_5_netPar2[2]}), .R_condition(rc[55]), .OUT(dalpha_L1_j_5[2]), .SIGN_out(SIGN_dalpha_L1_j_5[2]));
SS_ADDSUB ADDSUB_dalpha_L1_2_6(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_6_netPar0[2], dalpha_L1_j_6_netPar1[2], dalpha_L1_j_6_netPar2[2] }), .SIGN({ SIGN_dalpha_L1_j_6_netPar0[2], SIGN_dalpha_L1_j_6_netPar1[2], SIGN_dalpha_L1_j_6_netPar2[2]}), .R_condition(rc[56]), .OUT(dalpha_L1_j_6[2]), .SIGN_out(SIGN_dalpha_L1_j_6[2]));
SS_ADDSUB ADDSUB_dalpha_L1_2_7(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_7_netPar0[2], dalpha_L1_j_7_netPar1[2], dalpha_L1_j_7_netPar2[2] }), .SIGN({ SIGN_dalpha_L1_j_7_netPar0[2], SIGN_dalpha_L1_j_7_netPar1[2], SIGN_dalpha_L1_j_7_netPar2[2]}), .R_condition(rc[57]), .OUT(dalpha_L1_j_7[2]), .SIGN_out(SIGN_dalpha_L1_j_7[2]));
SS_ADDSUB ADDSUB_dalpha_L1_2_8(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_8_netPar0[2], dalpha_L1_j_8_netPar1[2], dalpha_L1_j_8_netPar2[2] }), .SIGN({ SIGN_dalpha_L1_j_8_netPar0[2], SIGN_dalpha_L1_j_8_netPar1[2], SIGN_dalpha_L1_j_8_netPar2[2]}), .R_condition(rc[58]), .OUT(dalpha_L1_j_8[2]), .SIGN_out(SIGN_dalpha_L1_j_8[2]));
SS_ADDSUB ADDSUB_dalpha_L1_2_9(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_9_netPar0[2], dalpha_L1_j_9_netPar1[2], dalpha_L1_j_9_netPar2[2] }), .SIGN({ SIGN_dalpha_L1_j_9_netPar0[2], SIGN_dalpha_L1_j_9_netPar1[2], SIGN_dalpha_L1_j_9_netPar2[2]}), .R_condition(rc[59]), .OUT(dalpha_L1_j_9[2]), .SIGN_out(SIGN_dalpha_L1_j_9[2]));
SS_ADDSUB ADDSUB_dalpha_L1_2_10(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_10_netPar0[2], dalpha_L1_j_10_netPar1[2], dalpha_L1_j_10_netPar2[2] }), .SIGN({ SIGN_dalpha_L1_j_10_netPar0[2], SIGN_dalpha_L1_j_10_netPar1[2], SIGN_dalpha_L1_j_10_netPar2[2]}), .R_condition(rc[60]), .OUT(dalpha_L1_j_10[2]), .SIGN_out(SIGN_dalpha_L1_j_10[2]));
SS_ADDSUB ADDSUB_dalpha_L1_2_11(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_11_netPar0[2], dalpha_L1_j_11_netPar1[2], dalpha_L1_j_11_netPar2[2] }), .SIGN({ SIGN_dalpha_L1_j_11_netPar0[2], SIGN_dalpha_L1_j_11_netPar1[2], SIGN_dalpha_L1_j_11_netPar2[2]}), .R_condition(rc[61]), .OUT(dalpha_L1_j_11[2]), .SIGN_out(SIGN_dalpha_L1_j_11[2]));
SS_ADDSUB ADDSUB_dalpha_L1_2_12(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_12_netPar0[2], dalpha_L1_j_12_netPar1[2], dalpha_L1_j_12_netPar2[2] }), .SIGN({ SIGN_dalpha_L1_j_12_netPar0[2], SIGN_dalpha_L1_j_12_netPar1[2], SIGN_dalpha_L1_j_12_netPar2[2]}), .R_condition(rc[62]), .OUT(dalpha_L1_j_12[2]), .SIGN_out(SIGN_dalpha_L1_j_12[2]));
SS_ADDSUB ADDSUB_dalpha_L1_2_13(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_13_netPar0[2], dalpha_L1_j_13_netPar1[2], dalpha_L1_j_13_netPar2[2] }), .SIGN({ SIGN_dalpha_L1_j_13_netPar0[2], SIGN_dalpha_L1_j_13_netPar1[2], SIGN_dalpha_L1_j_13_netPar2[2]}), .R_condition(rc[63]), .OUT(dalpha_L1_j_13[2]), .SIGN_out(SIGN_dalpha_L1_j_13[2]));
SS_ADDSUB ADDSUB_dalpha_L1_2_14(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_14_netPar0[2], dalpha_L1_j_14_netPar1[2], dalpha_L1_j_14_netPar2[2] }), .SIGN({ SIGN_dalpha_L1_j_14_netPar0[2], SIGN_dalpha_L1_j_14_netPar1[2], SIGN_dalpha_L1_j_14_netPar2[2]}), .R_condition(rc[64]), .OUT(dalpha_L1_j_14[2]), .SIGN_out(SIGN_dalpha_L1_j_14[2]));
SS_ADDSUB ADDSUB_dalpha_L1_2_15(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_15_netPar0[2], dalpha_L1_j_15_netPar1[2], dalpha_L1_j_15_netPar2[2] }), .SIGN({ SIGN_dalpha_L1_j_15_netPar0[2], SIGN_dalpha_L1_j_15_netPar1[2], SIGN_dalpha_L1_j_15_netPar2[2]}), .R_condition(rc[65]), .OUT(dalpha_L1_j_15[2]), .SIGN_out(SIGN_dalpha_L1_j_15[2]));
SS_ADDSUB ADDSUB_dalpha_L1_2_16(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_16_netPar0[2], dalpha_L1_j_16_netPar1[2], dalpha_L1_j_16_netPar2[2] }), .SIGN({ SIGN_dalpha_L1_j_16_netPar0[2], SIGN_dalpha_L1_j_16_netPar1[2], SIGN_dalpha_L1_j_16_netPar2[2]}), .R_condition(rc[66]), .OUT(dalpha_L1_j_16[2]), .SIGN_out(SIGN_dalpha_L1_j_16[2]));
SS_ADDSUB ADDSUB_dalpha_L1_2_17(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_17_netPar0[2], dalpha_L1_j_17_netPar1[2], dalpha_L1_j_17_netPar2[2] }), .SIGN({ SIGN_dalpha_L1_j_17_netPar0[2], SIGN_dalpha_L1_j_17_netPar1[2], SIGN_dalpha_L1_j_17_netPar2[2]}), .R_condition(rc[67]), .OUT(dalpha_L1_j_17[2]), .SIGN_out(SIGN_dalpha_L1_j_17[2]));
SS_ADDSUB ADDSUB_dalpha_L1_2_18(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_18_netPar0[2], dalpha_L1_j_18_netPar1[2], dalpha_L1_j_18_netPar2[2] }), .SIGN({ SIGN_dalpha_L1_j_18_netPar0[2], SIGN_dalpha_L1_j_18_netPar1[2], SIGN_dalpha_L1_j_18_netPar2[2]}), .R_condition(rc[68]), .OUT(dalpha_L1_j_18[2]), .SIGN_out(SIGN_dalpha_L1_j_18[2]));
SS_ADDSUB ADDSUB_dalpha_L1_2_19(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_19_netPar0[2], dalpha_L1_j_19_netPar1[2], dalpha_L1_j_19_netPar2[2] }), .SIGN({ SIGN_dalpha_L1_j_19_netPar0[2], SIGN_dalpha_L1_j_19_netPar1[2], SIGN_dalpha_L1_j_19_netPar2[2]}), .R_condition(rc[69]), .OUT(dalpha_L1_j_19[2]), .SIGN_out(SIGN_dalpha_L1_j_19[2]));
SS_ADDSUB ADDSUB_dalpha_L1_2_20(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_20_netPar0[2], dalpha_L1_j_20_netPar1[2], dalpha_L1_j_20_netPar2[2] }), .SIGN({ SIGN_dalpha_L1_j_20_netPar0[2], SIGN_dalpha_L1_j_20_netPar1[2], SIGN_dalpha_L1_j_20_netPar2[2]}), .R_condition(rc[70]), .OUT(dalpha_L1_j_20[2]), .SIGN_out(SIGN_dalpha_L1_j_20[2]));
SS_ADDSUB ADDSUB_dalpha_L1_2_21(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_21_netPar0[2], dalpha_L1_j_21_netPar1[2], dalpha_L1_j_21_netPar2[2] }), .SIGN({ SIGN_dalpha_L1_j_21_netPar0[2], SIGN_dalpha_L1_j_21_netPar1[2], SIGN_dalpha_L1_j_21_netPar2[2]}), .R_condition(rc[71]), .OUT(dalpha_L1_j_21[2]), .SIGN_out(SIGN_dalpha_L1_j_21[2]));
SS_ADDSUB ADDSUB_dalpha_L1_2_22(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_22_netPar0[2], dalpha_L1_j_22_netPar1[2], dalpha_L1_j_22_netPar2[2] }), .SIGN({ SIGN_dalpha_L1_j_22_netPar0[2], SIGN_dalpha_L1_j_22_netPar1[2], SIGN_dalpha_L1_j_22_netPar2[2]}), .R_condition(rc[72]), .OUT(dalpha_L1_j_22[2]), .SIGN_out(SIGN_dalpha_L1_j_22[2]));
SS_ADDSUB ADDSUB_dalpha_L1_2_23(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_23_netPar0[2], dalpha_L1_j_23_netPar1[2], dalpha_L1_j_23_netPar2[2] }), .SIGN({ SIGN_dalpha_L1_j_23_netPar0[2], SIGN_dalpha_L1_j_23_netPar1[2], SIGN_dalpha_L1_j_23_netPar2[2]}), .R_condition(rc[73]), .OUT(dalpha_L1_j_23[2]), .SIGN_out(SIGN_dalpha_L1_j_23[2]));
SS_ADDSUB ADDSUB_dalpha_L1_2_24(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_24_netPar0[2], dalpha_L1_j_24_netPar1[2], dalpha_L1_j_24_netPar2[2] }), .SIGN({ SIGN_dalpha_L1_j_24_netPar0[2], SIGN_dalpha_L1_j_24_netPar1[2], SIGN_dalpha_L1_j_24_netPar2[2]}), .R_condition(rc[74]), .OUT(dalpha_L1_j_24[2]), .SIGN_out(SIGN_dalpha_L1_j_24[2]));
SS_ADDSUB ADDSUB_dalpha_L1_3_0(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_0_netPar0[3], dalpha_L1_j_0_netPar1[3], dalpha_L1_j_0_netPar2[3] }), .SIGN({ SIGN_dalpha_L1_j_0_netPar0[3], SIGN_dalpha_L1_j_0_netPar1[3], SIGN_dalpha_L1_j_0_netPar2[3]}), .R_condition(rc[75]), .OUT(dalpha_L1_j_0[3]), .SIGN_out(SIGN_dalpha_L1_j_0[3]));
SS_ADDSUB ADDSUB_dalpha_L1_3_1(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_1_netPar0[3], dalpha_L1_j_1_netPar1[3], dalpha_L1_j_1_netPar2[3] }), .SIGN({ SIGN_dalpha_L1_j_1_netPar0[3], SIGN_dalpha_L1_j_1_netPar1[3], SIGN_dalpha_L1_j_1_netPar2[3]}), .R_condition(rc[76]), .OUT(dalpha_L1_j_1[3]), .SIGN_out(SIGN_dalpha_L1_j_1[3]));
SS_ADDSUB ADDSUB_dalpha_L1_3_2(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_2_netPar0[3], dalpha_L1_j_2_netPar1[3], dalpha_L1_j_2_netPar2[3] }), .SIGN({ SIGN_dalpha_L1_j_2_netPar0[3], SIGN_dalpha_L1_j_2_netPar1[3], SIGN_dalpha_L1_j_2_netPar2[3]}), .R_condition(rc[77]), .OUT(dalpha_L1_j_2[3]), .SIGN_out(SIGN_dalpha_L1_j_2[3]));
SS_ADDSUB ADDSUB_dalpha_L1_3_3(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_3_netPar0[3], dalpha_L1_j_3_netPar1[3], dalpha_L1_j_3_netPar2[3] }), .SIGN({ SIGN_dalpha_L1_j_3_netPar0[3], SIGN_dalpha_L1_j_3_netPar1[3], SIGN_dalpha_L1_j_3_netPar2[3]}), .R_condition(rc[78]), .OUT(dalpha_L1_j_3[3]), .SIGN_out(SIGN_dalpha_L1_j_3[3]));
SS_ADDSUB ADDSUB_dalpha_L1_3_4(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_4_netPar0[3], dalpha_L1_j_4_netPar1[3], dalpha_L1_j_4_netPar2[3] }), .SIGN({ SIGN_dalpha_L1_j_4_netPar0[3], SIGN_dalpha_L1_j_4_netPar1[3], SIGN_dalpha_L1_j_4_netPar2[3]}), .R_condition(rc[79]), .OUT(dalpha_L1_j_4[3]), .SIGN_out(SIGN_dalpha_L1_j_4[3]));
SS_ADDSUB ADDSUB_dalpha_L1_3_5(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_5_netPar0[3], dalpha_L1_j_5_netPar1[3], dalpha_L1_j_5_netPar2[3] }), .SIGN({ SIGN_dalpha_L1_j_5_netPar0[3], SIGN_dalpha_L1_j_5_netPar1[3], SIGN_dalpha_L1_j_5_netPar2[3]}), .R_condition(rc[80]), .OUT(dalpha_L1_j_5[3]), .SIGN_out(SIGN_dalpha_L1_j_5[3]));
SS_ADDSUB ADDSUB_dalpha_L1_3_6(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_6_netPar0[3], dalpha_L1_j_6_netPar1[3], dalpha_L1_j_6_netPar2[3] }), .SIGN({ SIGN_dalpha_L1_j_6_netPar0[3], SIGN_dalpha_L1_j_6_netPar1[3], SIGN_dalpha_L1_j_6_netPar2[3]}), .R_condition(rc[81]), .OUT(dalpha_L1_j_6[3]), .SIGN_out(SIGN_dalpha_L1_j_6[3]));
SS_ADDSUB ADDSUB_dalpha_L1_3_7(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_7_netPar0[3], dalpha_L1_j_7_netPar1[3], dalpha_L1_j_7_netPar2[3] }), .SIGN({ SIGN_dalpha_L1_j_7_netPar0[3], SIGN_dalpha_L1_j_7_netPar1[3], SIGN_dalpha_L1_j_7_netPar2[3]}), .R_condition(rc[82]), .OUT(dalpha_L1_j_7[3]), .SIGN_out(SIGN_dalpha_L1_j_7[3]));
SS_ADDSUB ADDSUB_dalpha_L1_3_8(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_8_netPar0[3], dalpha_L1_j_8_netPar1[3], dalpha_L1_j_8_netPar2[3] }), .SIGN({ SIGN_dalpha_L1_j_8_netPar0[3], SIGN_dalpha_L1_j_8_netPar1[3], SIGN_dalpha_L1_j_8_netPar2[3]}), .R_condition(rc[83]), .OUT(dalpha_L1_j_8[3]), .SIGN_out(SIGN_dalpha_L1_j_8[3]));
SS_ADDSUB ADDSUB_dalpha_L1_3_9(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_9_netPar0[3], dalpha_L1_j_9_netPar1[3], dalpha_L1_j_9_netPar2[3] }), .SIGN({ SIGN_dalpha_L1_j_9_netPar0[3], SIGN_dalpha_L1_j_9_netPar1[3], SIGN_dalpha_L1_j_9_netPar2[3]}), .R_condition(rc[84]), .OUT(dalpha_L1_j_9[3]), .SIGN_out(SIGN_dalpha_L1_j_9[3]));
SS_ADDSUB ADDSUB_dalpha_L1_3_10(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_10_netPar0[3], dalpha_L1_j_10_netPar1[3], dalpha_L1_j_10_netPar2[3] }), .SIGN({ SIGN_dalpha_L1_j_10_netPar0[3], SIGN_dalpha_L1_j_10_netPar1[3], SIGN_dalpha_L1_j_10_netPar2[3]}), .R_condition(rc[85]), .OUT(dalpha_L1_j_10[3]), .SIGN_out(SIGN_dalpha_L1_j_10[3]));
SS_ADDSUB ADDSUB_dalpha_L1_3_11(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_11_netPar0[3], dalpha_L1_j_11_netPar1[3], dalpha_L1_j_11_netPar2[3] }), .SIGN({ SIGN_dalpha_L1_j_11_netPar0[3], SIGN_dalpha_L1_j_11_netPar1[3], SIGN_dalpha_L1_j_11_netPar2[3]}), .R_condition(rc[86]), .OUT(dalpha_L1_j_11[3]), .SIGN_out(SIGN_dalpha_L1_j_11[3]));
SS_ADDSUB ADDSUB_dalpha_L1_3_12(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_12_netPar0[3], dalpha_L1_j_12_netPar1[3], dalpha_L1_j_12_netPar2[3] }), .SIGN({ SIGN_dalpha_L1_j_12_netPar0[3], SIGN_dalpha_L1_j_12_netPar1[3], SIGN_dalpha_L1_j_12_netPar2[3]}), .R_condition(rc[87]), .OUT(dalpha_L1_j_12[3]), .SIGN_out(SIGN_dalpha_L1_j_12[3]));
SS_ADDSUB ADDSUB_dalpha_L1_3_13(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_13_netPar0[3], dalpha_L1_j_13_netPar1[3], dalpha_L1_j_13_netPar2[3] }), .SIGN({ SIGN_dalpha_L1_j_13_netPar0[3], SIGN_dalpha_L1_j_13_netPar1[3], SIGN_dalpha_L1_j_13_netPar2[3]}), .R_condition(rc[88]), .OUT(dalpha_L1_j_13[3]), .SIGN_out(SIGN_dalpha_L1_j_13[3]));
SS_ADDSUB ADDSUB_dalpha_L1_3_14(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_14_netPar0[3], dalpha_L1_j_14_netPar1[3], dalpha_L1_j_14_netPar2[3] }), .SIGN({ SIGN_dalpha_L1_j_14_netPar0[3], SIGN_dalpha_L1_j_14_netPar1[3], SIGN_dalpha_L1_j_14_netPar2[3]}), .R_condition(rc[89]), .OUT(dalpha_L1_j_14[3]), .SIGN_out(SIGN_dalpha_L1_j_14[3]));
SS_ADDSUB ADDSUB_dalpha_L1_3_15(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_15_netPar0[3], dalpha_L1_j_15_netPar1[3], dalpha_L1_j_15_netPar2[3] }), .SIGN({ SIGN_dalpha_L1_j_15_netPar0[3], SIGN_dalpha_L1_j_15_netPar1[3], SIGN_dalpha_L1_j_15_netPar2[3]}), .R_condition(rc[90]), .OUT(dalpha_L1_j_15[3]), .SIGN_out(SIGN_dalpha_L1_j_15[3]));
SS_ADDSUB ADDSUB_dalpha_L1_3_16(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_16_netPar0[3], dalpha_L1_j_16_netPar1[3], dalpha_L1_j_16_netPar2[3] }), .SIGN({ SIGN_dalpha_L1_j_16_netPar0[3], SIGN_dalpha_L1_j_16_netPar1[3], SIGN_dalpha_L1_j_16_netPar2[3]}), .R_condition(rc[91]), .OUT(dalpha_L1_j_16[3]), .SIGN_out(SIGN_dalpha_L1_j_16[3]));
SS_ADDSUB ADDSUB_dalpha_L1_3_17(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_17_netPar0[3], dalpha_L1_j_17_netPar1[3], dalpha_L1_j_17_netPar2[3] }), .SIGN({ SIGN_dalpha_L1_j_17_netPar0[3], SIGN_dalpha_L1_j_17_netPar1[3], SIGN_dalpha_L1_j_17_netPar2[3]}), .R_condition(rc[92]), .OUT(dalpha_L1_j_17[3]), .SIGN_out(SIGN_dalpha_L1_j_17[3]));
SS_ADDSUB ADDSUB_dalpha_L1_3_18(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_18_netPar0[3], dalpha_L1_j_18_netPar1[3], dalpha_L1_j_18_netPar2[3] }), .SIGN({ SIGN_dalpha_L1_j_18_netPar0[3], SIGN_dalpha_L1_j_18_netPar1[3], SIGN_dalpha_L1_j_18_netPar2[3]}), .R_condition(rc[93]), .OUT(dalpha_L1_j_18[3]), .SIGN_out(SIGN_dalpha_L1_j_18[3]));
SS_ADDSUB ADDSUB_dalpha_L1_3_19(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_19_netPar0[3], dalpha_L1_j_19_netPar1[3], dalpha_L1_j_19_netPar2[3] }), .SIGN({ SIGN_dalpha_L1_j_19_netPar0[3], SIGN_dalpha_L1_j_19_netPar1[3], SIGN_dalpha_L1_j_19_netPar2[3]}), .R_condition(rc[94]), .OUT(dalpha_L1_j_19[3]), .SIGN_out(SIGN_dalpha_L1_j_19[3]));
SS_ADDSUB ADDSUB_dalpha_L1_3_20(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_20_netPar0[3], dalpha_L1_j_20_netPar1[3], dalpha_L1_j_20_netPar2[3] }), .SIGN({ SIGN_dalpha_L1_j_20_netPar0[3], SIGN_dalpha_L1_j_20_netPar1[3], SIGN_dalpha_L1_j_20_netPar2[3]}), .R_condition(rc[95]), .OUT(dalpha_L1_j_20[3]), .SIGN_out(SIGN_dalpha_L1_j_20[3]));
SS_ADDSUB ADDSUB_dalpha_L1_3_21(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_21_netPar0[3], dalpha_L1_j_21_netPar1[3], dalpha_L1_j_21_netPar2[3] }), .SIGN({ SIGN_dalpha_L1_j_21_netPar0[3], SIGN_dalpha_L1_j_21_netPar1[3], SIGN_dalpha_L1_j_21_netPar2[3]}), .R_condition(rc[96]), .OUT(dalpha_L1_j_21[3]), .SIGN_out(SIGN_dalpha_L1_j_21[3]));
SS_ADDSUB ADDSUB_dalpha_L1_3_22(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_22_netPar0[3], dalpha_L1_j_22_netPar1[3], dalpha_L1_j_22_netPar2[3] }), .SIGN({ SIGN_dalpha_L1_j_22_netPar0[3], SIGN_dalpha_L1_j_22_netPar1[3], SIGN_dalpha_L1_j_22_netPar2[3]}), .R_condition(rc[97]), .OUT(dalpha_L1_j_22[3]), .SIGN_out(SIGN_dalpha_L1_j_22[3]));
SS_ADDSUB ADDSUB_dalpha_L1_3_23(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_23_netPar0[3], dalpha_L1_j_23_netPar1[3], dalpha_L1_j_23_netPar2[3] }), .SIGN({ SIGN_dalpha_L1_j_23_netPar0[3], SIGN_dalpha_L1_j_23_netPar1[3], SIGN_dalpha_L1_j_23_netPar2[3]}), .R_condition(rc[98]), .OUT(dalpha_L1_j_23[3]), .SIGN_out(SIGN_dalpha_L1_j_23[3]));
SS_ADDSUB ADDSUB_dalpha_L1_3_24(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_24_netPar0[3], dalpha_L1_j_24_netPar1[3], dalpha_L1_j_24_netPar2[3] }), .SIGN({ SIGN_dalpha_L1_j_24_netPar0[3], SIGN_dalpha_L1_j_24_netPar1[3], SIGN_dalpha_L1_j_24_netPar2[3]}), .R_condition(rc[99]), .OUT(dalpha_L1_j_24[3]), .SIGN_out(SIGN_dalpha_L1_j_24[3]));
SS_ADDSUB ADDSUB_dalpha_L1_4_0(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_0_netPar0[4], dalpha_L1_j_0_netPar1[4], dalpha_L1_j_0_netPar2[4] }), .SIGN({ SIGN_dalpha_L1_j_0_netPar0[4], SIGN_dalpha_L1_j_0_netPar1[4], SIGN_dalpha_L1_j_0_netPar2[4]}), .R_condition(rc[100]), .OUT(dalpha_L1_j_0[4]), .SIGN_out(SIGN_dalpha_L1_j_0[4]));
SS_ADDSUB ADDSUB_dalpha_L1_4_1(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_1_netPar0[4], dalpha_L1_j_1_netPar1[4], dalpha_L1_j_1_netPar2[4] }), .SIGN({ SIGN_dalpha_L1_j_1_netPar0[4], SIGN_dalpha_L1_j_1_netPar1[4], SIGN_dalpha_L1_j_1_netPar2[4]}), .R_condition(rc[101]), .OUT(dalpha_L1_j_1[4]), .SIGN_out(SIGN_dalpha_L1_j_1[4]));
SS_ADDSUB ADDSUB_dalpha_L1_4_2(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_2_netPar0[4], dalpha_L1_j_2_netPar1[4], dalpha_L1_j_2_netPar2[4] }), .SIGN({ SIGN_dalpha_L1_j_2_netPar0[4], SIGN_dalpha_L1_j_2_netPar1[4], SIGN_dalpha_L1_j_2_netPar2[4]}), .R_condition(rc[102]), .OUT(dalpha_L1_j_2[4]), .SIGN_out(SIGN_dalpha_L1_j_2[4]));
SS_ADDSUB ADDSUB_dalpha_L1_4_3(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_3_netPar0[4], dalpha_L1_j_3_netPar1[4], dalpha_L1_j_3_netPar2[4] }), .SIGN({ SIGN_dalpha_L1_j_3_netPar0[4], SIGN_dalpha_L1_j_3_netPar1[4], SIGN_dalpha_L1_j_3_netPar2[4]}), .R_condition(rc[103]), .OUT(dalpha_L1_j_3[4]), .SIGN_out(SIGN_dalpha_L1_j_3[4]));
SS_ADDSUB ADDSUB_dalpha_L1_4_4(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_4_netPar0[4], dalpha_L1_j_4_netPar1[4], dalpha_L1_j_4_netPar2[4] }), .SIGN({ SIGN_dalpha_L1_j_4_netPar0[4], SIGN_dalpha_L1_j_4_netPar1[4], SIGN_dalpha_L1_j_4_netPar2[4]}), .R_condition(rc[104]), .OUT(dalpha_L1_j_4[4]), .SIGN_out(SIGN_dalpha_L1_j_4[4]));
SS_ADDSUB ADDSUB_dalpha_L1_4_5(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_5_netPar0[4], dalpha_L1_j_5_netPar1[4], dalpha_L1_j_5_netPar2[4] }), .SIGN({ SIGN_dalpha_L1_j_5_netPar0[4], SIGN_dalpha_L1_j_5_netPar1[4], SIGN_dalpha_L1_j_5_netPar2[4]}), .R_condition(rc[105]), .OUT(dalpha_L1_j_5[4]), .SIGN_out(SIGN_dalpha_L1_j_5[4]));
SS_ADDSUB ADDSUB_dalpha_L1_4_6(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_6_netPar0[4], dalpha_L1_j_6_netPar1[4], dalpha_L1_j_6_netPar2[4] }), .SIGN({ SIGN_dalpha_L1_j_6_netPar0[4], SIGN_dalpha_L1_j_6_netPar1[4], SIGN_dalpha_L1_j_6_netPar2[4]}), .R_condition(rc[106]), .OUT(dalpha_L1_j_6[4]), .SIGN_out(SIGN_dalpha_L1_j_6[4]));
SS_ADDSUB ADDSUB_dalpha_L1_4_7(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_7_netPar0[4], dalpha_L1_j_7_netPar1[4], dalpha_L1_j_7_netPar2[4] }), .SIGN({ SIGN_dalpha_L1_j_7_netPar0[4], SIGN_dalpha_L1_j_7_netPar1[4], SIGN_dalpha_L1_j_7_netPar2[4]}), .R_condition(rc[107]), .OUT(dalpha_L1_j_7[4]), .SIGN_out(SIGN_dalpha_L1_j_7[4]));
SS_ADDSUB ADDSUB_dalpha_L1_4_8(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_8_netPar0[4], dalpha_L1_j_8_netPar1[4], dalpha_L1_j_8_netPar2[4] }), .SIGN({ SIGN_dalpha_L1_j_8_netPar0[4], SIGN_dalpha_L1_j_8_netPar1[4], SIGN_dalpha_L1_j_8_netPar2[4]}), .R_condition(rc[108]), .OUT(dalpha_L1_j_8[4]), .SIGN_out(SIGN_dalpha_L1_j_8[4]));
SS_ADDSUB ADDSUB_dalpha_L1_4_9(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_9_netPar0[4], dalpha_L1_j_9_netPar1[4], dalpha_L1_j_9_netPar2[4] }), .SIGN({ SIGN_dalpha_L1_j_9_netPar0[4], SIGN_dalpha_L1_j_9_netPar1[4], SIGN_dalpha_L1_j_9_netPar2[4]}), .R_condition(rc[109]), .OUT(dalpha_L1_j_9[4]), .SIGN_out(SIGN_dalpha_L1_j_9[4]));
SS_ADDSUB ADDSUB_dalpha_L1_4_10(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_10_netPar0[4], dalpha_L1_j_10_netPar1[4], dalpha_L1_j_10_netPar2[4] }), .SIGN({ SIGN_dalpha_L1_j_10_netPar0[4], SIGN_dalpha_L1_j_10_netPar1[4], SIGN_dalpha_L1_j_10_netPar2[4]}), .R_condition(rc[110]), .OUT(dalpha_L1_j_10[4]), .SIGN_out(SIGN_dalpha_L1_j_10[4]));
SS_ADDSUB ADDSUB_dalpha_L1_4_11(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_11_netPar0[4], dalpha_L1_j_11_netPar1[4], dalpha_L1_j_11_netPar2[4] }), .SIGN({ SIGN_dalpha_L1_j_11_netPar0[4], SIGN_dalpha_L1_j_11_netPar1[4], SIGN_dalpha_L1_j_11_netPar2[4]}), .R_condition(rc[111]), .OUT(dalpha_L1_j_11[4]), .SIGN_out(SIGN_dalpha_L1_j_11[4]));
SS_ADDSUB ADDSUB_dalpha_L1_4_12(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_12_netPar0[4], dalpha_L1_j_12_netPar1[4], dalpha_L1_j_12_netPar2[4] }), .SIGN({ SIGN_dalpha_L1_j_12_netPar0[4], SIGN_dalpha_L1_j_12_netPar1[4], SIGN_dalpha_L1_j_12_netPar2[4]}), .R_condition(rc[112]), .OUT(dalpha_L1_j_12[4]), .SIGN_out(SIGN_dalpha_L1_j_12[4]));
SS_ADDSUB ADDSUB_dalpha_L1_4_13(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_13_netPar0[4], dalpha_L1_j_13_netPar1[4], dalpha_L1_j_13_netPar2[4] }), .SIGN({ SIGN_dalpha_L1_j_13_netPar0[4], SIGN_dalpha_L1_j_13_netPar1[4], SIGN_dalpha_L1_j_13_netPar2[4]}), .R_condition(rc[113]), .OUT(dalpha_L1_j_13[4]), .SIGN_out(SIGN_dalpha_L1_j_13[4]));
SS_ADDSUB ADDSUB_dalpha_L1_4_14(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_14_netPar0[4], dalpha_L1_j_14_netPar1[4], dalpha_L1_j_14_netPar2[4] }), .SIGN({ SIGN_dalpha_L1_j_14_netPar0[4], SIGN_dalpha_L1_j_14_netPar1[4], SIGN_dalpha_L1_j_14_netPar2[4]}), .R_condition(rc[114]), .OUT(dalpha_L1_j_14[4]), .SIGN_out(SIGN_dalpha_L1_j_14[4]));
SS_ADDSUB ADDSUB_dalpha_L1_4_15(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_15_netPar0[4], dalpha_L1_j_15_netPar1[4], dalpha_L1_j_15_netPar2[4] }), .SIGN({ SIGN_dalpha_L1_j_15_netPar0[4], SIGN_dalpha_L1_j_15_netPar1[4], SIGN_dalpha_L1_j_15_netPar2[4]}), .R_condition(rc[115]), .OUT(dalpha_L1_j_15[4]), .SIGN_out(SIGN_dalpha_L1_j_15[4]));
SS_ADDSUB ADDSUB_dalpha_L1_4_16(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_16_netPar0[4], dalpha_L1_j_16_netPar1[4], dalpha_L1_j_16_netPar2[4] }), .SIGN({ SIGN_dalpha_L1_j_16_netPar0[4], SIGN_dalpha_L1_j_16_netPar1[4], SIGN_dalpha_L1_j_16_netPar2[4]}), .R_condition(rc[116]), .OUT(dalpha_L1_j_16[4]), .SIGN_out(SIGN_dalpha_L1_j_16[4]));
SS_ADDSUB ADDSUB_dalpha_L1_4_17(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_17_netPar0[4], dalpha_L1_j_17_netPar1[4], dalpha_L1_j_17_netPar2[4] }), .SIGN({ SIGN_dalpha_L1_j_17_netPar0[4], SIGN_dalpha_L1_j_17_netPar1[4], SIGN_dalpha_L1_j_17_netPar2[4]}), .R_condition(rc[117]), .OUT(dalpha_L1_j_17[4]), .SIGN_out(SIGN_dalpha_L1_j_17[4]));
SS_ADDSUB ADDSUB_dalpha_L1_4_18(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_18_netPar0[4], dalpha_L1_j_18_netPar1[4], dalpha_L1_j_18_netPar2[4] }), .SIGN({ SIGN_dalpha_L1_j_18_netPar0[4], SIGN_dalpha_L1_j_18_netPar1[4], SIGN_dalpha_L1_j_18_netPar2[4]}), .R_condition(rc[118]), .OUT(dalpha_L1_j_18[4]), .SIGN_out(SIGN_dalpha_L1_j_18[4]));
SS_ADDSUB ADDSUB_dalpha_L1_4_19(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_19_netPar0[4], dalpha_L1_j_19_netPar1[4], dalpha_L1_j_19_netPar2[4] }), .SIGN({ SIGN_dalpha_L1_j_19_netPar0[4], SIGN_dalpha_L1_j_19_netPar1[4], SIGN_dalpha_L1_j_19_netPar2[4]}), .R_condition(rc[119]), .OUT(dalpha_L1_j_19[4]), .SIGN_out(SIGN_dalpha_L1_j_19[4]));
SS_ADDSUB ADDSUB_dalpha_L1_4_20(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_20_netPar0[4], dalpha_L1_j_20_netPar1[4], dalpha_L1_j_20_netPar2[4] }), .SIGN({ SIGN_dalpha_L1_j_20_netPar0[4], SIGN_dalpha_L1_j_20_netPar1[4], SIGN_dalpha_L1_j_20_netPar2[4]}), .R_condition(rc[120]), .OUT(dalpha_L1_j_20[4]), .SIGN_out(SIGN_dalpha_L1_j_20[4]));
SS_ADDSUB ADDSUB_dalpha_L1_4_21(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_21_netPar0[4], dalpha_L1_j_21_netPar1[4], dalpha_L1_j_21_netPar2[4] }), .SIGN({ SIGN_dalpha_L1_j_21_netPar0[4], SIGN_dalpha_L1_j_21_netPar1[4], SIGN_dalpha_L1_j_21_netPar2[4]}), .R_condition(rc[121]), .OUT(dalpha_L1_j_21[4]), .SIGN_out(SIGN_dalpha_L1_j_21[4]));
SS_ADDSUB ADDSUB_dalpha_L1_4_22(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_22_netPar0[4], dalpha_L1_j_22_netPar1[4], dalpha_L1_j_22_netPar2[4] }), .SIGN({ SIGN_dalpha_L1_j_22_netPar0[4], SIGN_dalpha_L1_j_22_netPar1[4], SIGN_dalpha_L1_j_22_netPar2[4]}), .R_condition(rc[122]), .OUT(dalpha_L1_j_22[4]), .SIGN_out(SIGN_dalpha_L1_j_22[4]));
SS_ADDSUB ADDSUB_dalpha_L1_4_23(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_23_netPar0[4], dalpha_L1_j_23_netPar1[4], dalpha_L1_j_23_netPar2[4] }), .SIGN({ SIGN_dalpha_L1_j_23_netPar0[4], SIGN_dalpha_L1_j_23_netPar1[4], SIGN_dalpha_L1_j_23_netPar2[4]}), .R_condition(rc[123]), .OUT(dalpha_L1_j_23[4]), .SIGN_out(SIGN_dalpha_L1_j_23[4]));
SS_ADDSUB ADDSUB_dalpha_L1_4_24(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L1_j_24_netPar0[4], dalpha_L1_j_24_netPar1[4], dalpha_L1_j_24_netPar2[4] }), .SIGN({ SIGN_dalpha_L1_j_24_netPar0[4], SIGN_dalpha_L1_j_24_netPar1[4], SIGN_dalpha_L1_j_24_netPar2[4]}), .R_condition(rc[124]), .OUT(dalpha_L1_j_24[4]), .SIGN_out(SIGN_dalpha_L1_j_24[4]));
defparam ADDSUB_dalpha_L1_0_0.N = 3;
defparam ADDSUB_dalpha_L1_0_1.N = 3;
defparam ADDSUB_dalpha_L1_0_2.N = 3;
defparam ADDSUB_dalpha_L1_0_3.N = 3;
defparam ADDSUB_dalpha_L1_0_4.N = 3;
defparam ADDSUB_dalpha_L1_0_5.N = 3;
defparam ADDSUB_dalpha_L1_0_6.N = 3;
defparam ADDSUB_dalpha_L1_0_7.N = 3;
defparam ADDSUB_dalpha_L1_0_8.N = 3;
defparam ADDSUB_dalpha_L1_0_9.N = 3;
defparam ADDSUB_dalpha_L1_0_10.N = 3;
defparam ADDSUB_dalpha_L1_0_11.N = 3;
defparam ADDSUB_dalpha_L1_0_12.N = 3;
defparam ADDSUB_dalpha_L1_0_13.N = 3;
defparam ADDSUB_dalpha_L1_0_14.N = 3;
defparam ADDSUB_dalpha_L1_0_15.N = 3;
defparam ADDSUB_dalpha_L1_0_16.N = 3;
defparam ADDSUB_dalpha_L1_0_17.N = 3;
defparam ADDSUB_dalpha_L1_0_18.N = 3;
defparam ADDSUB_dalpha_L1_0_19.N = 3;
defparam ADDSUB_dalpha_L1_0_20.N = 3;
defparam ADDSUB_dalpha_L1_0_21.N = 3;
defparam ADDSUB_dalpha_L1_0_22.N = 3;
defparam ADDSUB_dalpha_L1_0_23.N = 3;
defparam ADDSUB_dalpha_L1_0_24.N = 3;
defparam ADDSUB_dalpha_L1_1_0.N = 3;
defparam ADDSUB_dalpha_L1_1_1.N = 3;
defparam ADDSUB_dalpha_L1_1_2.N = 3;
defparam ADDSUB_dalpha_L1_1_3.N = 3;
defparam ADDSUB_dalpha_L1_1_4.N = 3;
defparam ADDSUB_dalpha_L1_1_5.N = 3;
defparam ADDSUB_dalpha_L1_1_6.N = 3;
defparam ADDSUB_dalpha_L1_1_7.N = 3;
defparam ADDSUB_dalpha_L1_1_8.N = 3;
defparam ADDSUB_dalpha_L1_1_9.N = 3;
defparam ADDSUB_dalpha_L1_1_10.N = 3;
defparam ADDSUB_dalpha_L1_1_11.N = 3;
defparam ADDSUB_dalpha_L1_1_12.N = 3;
defparam ADDSUB_dalpha_L1_1_13.N = 3;
defparam ADDSUB_dalpha_L1_1_14.N = 3;
defparam ADDSUB_dalpha_L1_1_15.N = 3;
defparam ADDSUB_dalpha_L1_1_16.N = 3;
defparam ADDSUB_dalpha_L1_1_17.N = 3;
defparam ADDSUB_dalpha_L1_1_18.N = 3;
defparam ADDSUB_dalpha_L1_1_19.N = 3;
defparam ADDSUB_dalpha_L1_1_20.N = 3;
defparam ADDSUB_dalpha_L1_1_21.N = 3;
defparam ADDSUB_dalpha_L1_1_22.N = 3;
defparam ADDSUB_dalpha_L1_1_23.N = 3;
defparam ADDSUB_dalpha_L1_1_24.N = 3;
defparam ADDSUB_dalpha_L1_2_0.N = 3;
defparam ADDSUB_dalpha_L1_2_1.N = 3;
defparam ADDSUB_dalpha_L1_2_2.N = 3;
defparam ADDSUB_dalpha_L1_2_3.N = 3;
defparam ADDSUB_dalpha_L1_2_4.N = 3;
defparam ADDSUB_dalpha_L1_2_5.N = 3;
defparam ADDSUB_dalpha_L1_2_6.N = 3;
defparam ADDSUB_dalpha_L1_2_7.N = 3;
defparam ADDSUB_dalpha_L1_2_8.N = 3;
defparam ADDSUB_dalpha_L1_2_9.N = 3;
defparam ADDSUB_dalpha_L1_2_10.N = 3;
defparam ADDSUB_dalpha_L1_2_11.N = 3;
defparam ADDSUB_dalpha_L1_2_12.N = 3;
defparam ADDSUB_dalpha_L1_2_13.N = 3;
defparam ADDSUB_dalpha_L1_2_14.N = 3;
defparam ADDSUB_dalpha_L1_2_15.N = 3;
defparam ADDSUB_dalpha_L1_2_16.N = 3;
defparam ADDSUB_dalpha_L1_2_17.N = 3;
defparam ADDSUB_dalpha_L1_2_18.N = 3;
defparam ADDSUB_dalpha_L1_2_19.N = 3;
defparam ADDSUB_dalpha_L1_2_20.N = 3;
defparam ADDSUB_dalpha_L1_2_21.N = 3;
defparam ADDSUB_dalpha_L1_2_22.N = 3;
defparam ADDSUB_dalpha_L1_2_23.N = 3;
defparam ADDSUB_dalpha_L1_2_24.N = 3;
defparam ADDSUB_dalpha_L1_3_0.N = 3;
defparam ADDSUB_dalpha_L1_3_1.N = 3;
defparam ADDSUB_dalpha_L1_3_2.N = 3;
defparam ADDSUB_dalpha_L1_3_3.N = 3;
defparam ADDSUB_dalpha_L1_3_4.N = 3;
defparam ADDSUB_dalpha_L1_3_5.N = 3;
defparam ADDSUB_dalpha_L1_3_6.N = 3;
defparam ADDSUB_dalpha_L1_3_7.N = 3;
defparam ADDSUB_dalpha_L1_3_8.N = 3;
defparam ADDSUB_dalpha_L1_3_9.N = 3;
defparam ADDSUB_dalpha_L1_3_10.N = 3;
defparam ADDSUB_dalpha_L1_3_11.N = 3;
defparam ADDSUB_dalpha_L1_3_12.N = 3;
defparam ADDSUB_dalpha_L1_3_13.N = 3;
defparam ADDSUB_dalpha_L1_3_14.N = 3;
defparam ADDSUB_dalpha_L1_3_15.N = 3;
defparam ADDSUB_dalpha_L1_3_16.N = 3;
defparam ADDSUB_dalpha_L1_3_17.N = 3;
defparam ADDSUB_dalpha_L1_3_18.N = 3;
defparam ADDSUB_dalpha_L1_3_19.N = 3;
defparam ADDSUB_dalpha_L1_3_20.N = 3;
defparam ADDSUB_dalpha_L1_3_21.N = 3;
defparam ADDSUB_dalpha_L1_3_22.N = 3;
defparam ADDSUB_dalpha_L1_3_23.N = 3;
defparam ADDSUB_dalpha_L1_3_24.N = 3;
defparam ADDSUB_dalpha_L1_4_0.N = 3;
defparam ADDSUB_dalpha_L1_4_1.N = 3;
defparam ADDSUB_dalpha_L1_4_2.N = 3;
defparam ADDSUB_dalpha_L1_4_3.N = 3;
defparam ADDSUB_dalpha_L1_4_4.N = 3;
defparam ADDSUB_dalpha_L1_4_5.N = 3;
defparam ADDSUB_dalpha_L1_4_6.N = 3;
defparam ADDSUB_dalpha_L1_4_7.N = 3;
defparam ADDSUB_dalpha_L1_4_8.N = 3;
defparam ADDSUB_dalpha_L1_4_9.N = 3;
defparam ADDSUB_dalpha_L1_4_10.N = 3;
defparam ADDSUB_dalpha_L1_4_11.N = 3;
defparam ADDSUB_dalpha_L1_4_12.N = 3;
defparam ADDSUB_dalpha_L1_4_13.N = 3;
defparam ADDSUB_dalpha_L1_4_14.N = 3;
defparam ADDSUB_dalpha_L1_4_15.N = 3;
defparam ADDSUB_dalpha_L1_4_16.N = 3;
defparam ADDSUB_dalpha_L1_4_17.N = 3;
defparam ADDSUB_dalpha_L1_4_18.N = 3;
defparam ADDSUB_dalpha_L1_4_19.N = 3;
defparam ADDSUB_dalpha_L1_4_20.N = 3;
defparam ADDSUB_dalpha_L1_4_21.N = 3;
defparam ADDSUB_dalpha_L1_4_22.N = 3;
defparam ADDSUB_dalpha_L1_4_23.N = 3;
defparam ADDSUB_dalpha_L1_4_24.N = 3;
defparam ADDSUB_dalpha_L1_0_0.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_0_1.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_0_2.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_0_3.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_0_4.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_0_5.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_0_6.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_0_7.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_0_8.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_0_9.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_0_10.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_0_11.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_0_12.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_0_13.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_0_14.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_0_15.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_0_16.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_0_17.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_0_18.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_0_19.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_0_20.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_0_21.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_0_22.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_0_23.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_0_24.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_1_0.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_1_1.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_1_2.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_1_3.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_1_4.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_1_5.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_1_6.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_1_7.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_1_8.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_1_9.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_1_10.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_1_11.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_1_12.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_1_13.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_1_14.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_1_15.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_1_16.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_1_17.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_1_18.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_1_19.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_1_20.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_1_21.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_1_22.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_1_23.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_1_24.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_2_0.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_2_1.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_2_2.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_2_3.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_2_4.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_2_5.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_2_6.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_2_7.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_2_8.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_2_9.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_2_10.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_2_11.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_2_12.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_2_13.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_2_14.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_2_15.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_2_16.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_2_17.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_2_18.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_2_19.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_2_20.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_2_21.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_2_22.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_2_23.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_2_24.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_3_0.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_3_1.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_3_2.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_3_3.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_3_4.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_3_5.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_3_6.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_3_7.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_3_8.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_3_9.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_3_10.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_3_11.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_3_12.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_3_13.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_3_14.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_3_15.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_3_16.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_3_17.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_3_18.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_3_19.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_3_20.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_3_21.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_3_22.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_3_23.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_3_24.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_4_0.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_4_1.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_4_2.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_4_3.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_4_4.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_4_5.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_4_6.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_4_7.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_4_8.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_4_9.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_4_10.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_4_11.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_4_12.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_4_13.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_4_14.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_4_15.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_4_16.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_4_17.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_4_18.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_4_19.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_4_20.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_4_21.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_4_22.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_4_23.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L1_4_24.DIFFCOUNTER_SIZE = 3;

SS_ADDSUB ADDSUB_dbeta_L1_0(.CLK(CLK), .INIT(INIT), .IN({ dbeta_L1_netPar0[0], dbeta_L1_netPar1[0], dbeta_L1_netPar2[0] }), .SIGN({ SIGN_dbeta_L1_netPar0[0], SIGN_dbeta_L1_netPar1[0], SIGN_dbeta_L1_netPar2[0]}), .R_condition(rc[125]), .OUT(dbeta_L1[0]), .SIGN_out(SIGN_dbeta_L1[0]));
SS_ADDSUB ADDSUB_dbeta_L1_1(.CLK(CLK), .INIT(INIT), .IN({ dbeta_L1_netPar0[1], dbeta_L1_netPar1[1], dbeta_L1_netPar2[1] }), .SIGN({ SIGN_dbeta_L1_netPar0[1], SIGN_dbeta_L1_netPar1[1], SIGN_dbeta_L1_netPar2[1]}), .R_condition(rc[126]), .OUT(dbeta_L1[1]), .SIGN_out(SIGN_dbeta_L1[1]));
SS_ADDSUB ADDSUB_dbeta_L1_2(.CLK(CLK), .INIT(INIT), .IN({ dbeta_L1_netPar0[2], dbeta_L1_netPar1[2], dbeta_L1_netPar2[2] }), .SIGN({ SIGN_dbeta_L1_netPar0[2], SIGN_dbeta_L1_netPar1[2], SIGN_dbeta_L1_netPar2[2]}), .R_condition(rc[127]), .OUT(dbeta_L1[2]), .SIGN_out(SIGN_dbeta_L1[2]));
SS_ADDSUB ADDSUB_dbeta_L1_3(.CLK(CLK), .INIT(INIT), .IN({ dbeta_L1_netPar0[3], dbeta_L1_netPar1[3], dbeta_L1_netPar2[3] }), .SIGN({ SIGN_dbeta_L1_netPar0[3], SIGN_dbeta_L1_netPar1[3], SIGN_dbeta_L1_netPar2[3]}), .R_condition(rc[128]), .OUT(dbeta_L1[3]), .SIGN_out(SIGN_dbeta_L1[3]));
SS_ADDSUB ADDSUB_dbeta_L1_4(.CLK(CLK), .INIT(INIT), .IN({ dbeta_L1_netPar0[4], dbeta_L1_netPar1[4], dbeta_L1_netPar2[4] }), .SIGN({ SIGN_dbeta_L1_netPar0[4], SIGN_dbeta_L1_netPar1[4], SIGN_dbeta_L1_netPar2[4]}), .R_condition(rc[129]), .OUT(dbeta_L1[4]), .SIGN_out(SIGN_dbeta_L1[4]));
SS_ADDSUB ADDSUB_dbeta_L1_5(.CLK(CLK), .INIT(INIT), .IN({ dbeta_L1_netPar0[5], dbeta_L1_netPar1[5], dbeta_L1_netPar2[5] }), .SIGN({ SIGN_dbeta_L1_netPar0[5], SIGN_dbeta_L1_netPar1[5], SIGN_dbeta_L1_netPar2[5]}), .R_condition(rc[130]), .OUT(dbeta_L1[5]), .SIGN_out(SIGN_dbeta_L1[5]));
SS_ADDSUB ADDSUB_dbeta_L1_6(.CLK(CLK), .INIT(INIT), .IN({ dbeta_L1_netPar0[6], dbeta_L1_netPar1[6], dbeta_L1_netPar2[6] }), .SIGN({ SIGN_dbeta_L1_netPar0[6], SIGN_dbeta_L1_netPar1[6], SIGN_dbeta_L1_netPar2[6]}), .R_condition(rc[131]), .OUT(dbeta_L1[6]), .SIGN_out(SIGN_dbeta_L1[6]));
SS_ADDSUB ADDSUB_dbeta_L1_7(.CLK(CLK), .INIT(INIT), .IN({ dbeta_L1_netPar0[7], dbeta_L1_netPar1[7], dbeta_L1_netPar2[7] }), .SIGN({ SIGN_dbeta_L1_netPar0[7], SIGN_dbeta_L1_netPar1[7], SIGN_dbeta_L1_netPar2[7]}), .R_condition(rc[132]), .OUT(dbeta_L1[7]), .SIGN_out(SIGN_dbeta_L1[7]));
SS_ADDSUB ADDSUB_dbeta_L1_8(.CLK(CLK), .INIT(INIT), .IN({ dbeta_L1_netPar0[8], dbeta_L1_netPar1[8], dbeta_L1_netPar2[8] }), .SIGN({ SIGN_dbeta_L1_netPar0[8], SIGN_dbeta_L1_netPar1[8], SIGN_dbeta_L1_netPar2[8]}), .R_condition(rc[133]), .OUT(dbeta_L1[8]), .SIGN_out(SIGN_dbeta_L1[8]));
SS_ADDSUB ADDSUB_dbeta_L1_9(.CLK(CLK), .INIT(INIT), .IN({ dbeta_L1_netPar0[9], dbeta_L1_netPar1[9], dbeta_L1_netPar2[9] }), .SIGN({ SIGN_dbeta_L1_netPar0[9], SIGN_dbeta_L1_netPar1[9], SIGN_dbeta_L1_netPar2[9]}), .R_condition(rc[134]), .OUT(dbeta_L1[9]), .SIGN_out(SIGN_dbeta_L1[9]));
SS_ADDSUB ADDSUB_dbeta_L1_10(.CLK(CLK), .INIT(INIT), .IN({ dbeta_L1_netPar0[10], dbeta_L1_netPar1[10], dbeta_L1_netPar2[10] }), .SIGN({ SIGN_dbeta_L1_netPar0[10], SIGN_dbeta_L1_netPar1[10], SIGN_dbeta_L1_netPar2[10]}), .R_condition(rc[135]), .OUT(dbeta_L1[10]), .SIGN_out(SIGN_dbeta_L1[10]));
SS_ADDSUB ADDSUB_dbeta_L1_11(.CLK(CLK), .INIT(INIT), .IN({ dbeta_L1_netPar0[11], dbeta_L1_netPar1[11], dbeta_L1_netPar2[11] }), .SIGN({ SIGN_dbeta_L1_netPar0[11], SIGN_dbeta_L1_netPar1[11], SIGN_dbeta_L1_netPar2[11]}), .R_condition(rc[136]), .OUT(dbeta_L1[11]), .SIGN_out(SIGN_dbeta_L1[11]));
SS_ADDSUB ADDSUB_dbeta_L1_12(.CLK(CLK), .INIT(INIT), .IN({ dbeta_L1_netPar0[12], dbeta_L1_netPar1[12], dbeta_L1_netPar2[12] }), .SIGN({ SIGN_dbeta_L1_netPar0[12], SIGN_dbeta_L1_netPar1[12], SIGN_dbeta_L1_netPar2[12]}), .R_condition(rc[137]), .OUT(dbeta_L1[12]), .SIGN_out(SIGN_dbeta_L1[12]));
SS_ADDSUB ADDSUB_dbeta_L1_13(.CLK(CLK), .INIT(INIT), .IN({ dbeta_L1_netPar0[13], dbeta_L1_netPar1[13], dbeta_L1_netPar2[13] }), .SIGN({ SIGN_dbeta_L1_netPar0[13], SIGN_dbeta_L1_netPar1[13], SIGN_dbeta_L1_netPar2[13]}), .R_condition(rc[138]), .OUT(dbeta_L1[13]), .SIGN_out(SIGN_dbeta_L1[13]));
SS_ADDSUB ADDSUB_dbeta_L1_14(.CLK(CLK), .INIT(INIT), .IN({ dbeta_L1_netPar0[14], dbeta_L1_netPar1[14], dbeta_L1_netPar2[14] }), .SIGN({ SIGN_dbeta_L1_netPar0[14], SIGN_dbeta_L1_netPar1[14], SIGN_dbeta_L1_netPar2[14]}), .R_condition(rc[139]), .OUT(dbeta_L1[14]), .SIGN_out(SIGN_dbeta_L1[14]));
SS_ADDSUB ADDSUB_dbeta_L1_15(.CLK(CLK), .INIT(INIT), .IN({ dbeta_L1_netPar0[15], dbeta_L1_netPar1[15], dbeta_L1_netPar2[15] }), .SIGN({ SIGN_dbeta_L1_netPar0[15], SIGN_dbeta_L1_netPar1[15], SIGN_dbeta_L1_netPar2[15]}), .R_condition(rc[140]), .OUT(dbeta_L1[15]), .SIGN_out(SIGN_dbeta_L1[15]));
SS_ADDSUB ADDSUB_dbeta_L1_16(.CLK(CLK), .INIT(INIT), .IN({ dbeta_L1_netPar0[16], dbeta_L1_netPar1[16], dbeta_L1_netPar2[16] }), .SIGN({ SIGN_dbeta_L1_netPar0[16], SIGN_dbeta_L1_netPar1[16], SIGN_dbeta_L1_netPar2[16]}), .R_condition(rc[141]), .OUT(dbeta_L1[16]), .SIGN_out(SIGN_dbeta_L1[16]));
SS_ADDSUB ADDSUB_dbeta_L1_17(.CLK(CLK), .INIT(INIT), .IN({ dbeta_L1_netPar0[17], dbeta_L1_netPar1[17], dbeta_L1_netPar2[17] }), .SIGN({ SIGN_dbeta_L1_netPar0[17], SIGN_dbeta_L1_netPar1[17], SIGN_dbeta_L1_netPar2[17]}), .R_condition(rc[142]), .OUT(dbeta_L1[17]), .SIGN_out(SIGN_dbeta_L1[17]));
SS_ADDSUB ADDSUB_dbeta_L1_18(.CLK(CLK), .INIT(INIT), .IN({ dbeta_L1_netPar0[18], dbeta_L1_netPar1[18], dbeta_L1_netPar2[18] }), .SIGN({ SIGN_dbeta_L1_netPar0[18], SIGN_dbeta_L1_netPar1[18], SIGN_dbeta_L1_netPar2[18]}), .R_condition(rc[143]), .OUT(dbeta_L1[18]), .SIGN_out(SIGN_dbeta_L1[18]));
SS_ADDSUB ADDSUB_dbeta_L1_19(.CLK(CLK), .INIT(INIT), .IN({ dbeta_L1_netPar0[19], dbeta_L1_netPar1[19], dbeta_L1_netPar2[19] }), .SIGN({ SIGN_dbeta_L1_netPar0[19], SIGN_dbeta_L1_netPar1[19], SIGN_dbeta_L1_netPar2[19]}), .R_condition(rc[144]), .OUT(dbeta_L1[19]), .SIGN_out(SIGN_dbeta_L1[19]));
SS_ADDSUB ADDSUB_dbeta_L1_20(.CLK(CLK), .INIT(INIT), .IN({ dbeta_L1_netPar0[20], dbeta_L1_netPar1[20], dbeta_L1_netPar2[20] }), .SIGN({ SIGN_dbeta_L1_netPar0[20], SIGN_dbeta_L1_netPar1[20], SIGN_dbeta_L1_netPar2[20]}), .R_condition(rc[145]), .OUT(dbeta_L1[20]), .SIGN_out(SIGN_dbeta_L1[20]));
SS_ADDSUB ADDSUB_dbeta_L1_21(.CLK(CLK), .INIT(INIT), .IN({ dbeta_L1_netPar0[21], dbeta_L1_netPar1[21], dbeta_L1_netPar2[21] }), .SIGN({ SIGN_dbeta_L1_netPar0[21], SIGN_dbeta_L1_netPar1[21], SIGN_dbeta_L1_netPar2[21]}), .R_condition(rc[146]), .OUT(dbeta_L1[21]), .SIGN_out(SIGN_dbeta_L1[21]));
SS_ADDSUB ADDSUB_dbeta_L1_22(.CLK(CLK), .INIT(INIT), .IN({ dbeta_L1_netPar0[22], dbeta_L1_netPar1[22], dbeta_L1_netPar2[22] }), .SIGN({ SIGN_dbeta_L1_netPar0[22], SIGN_dbeta_L1_netPar1[22], SIGN_dbeta_L1_netPar2[22]}), .R_condition(rc[147]), .OUT(dbeta_L1[22]), .SIGN_out(SIGN_dbeta_L1[22]));
SS_ADDSUB ADDSUB_dbeta_L1_23(.CLK(CLK), .INIT(INIT), .IN({ dbeta_L1_netPar0[23], dbeta_L1_netPar1[23], dbeta_L1_netPar2[23] }), .SIGN({ SIGN_dbeta_L1_netPar0[23], SIGN_dbeta_L1_netPar1[23], SIGN_dbeta_L1_netPar2[23]}), .R_condition(rc[148]), .OUT(dbeta_L1[23]), .SIGN_out(SIGN_dbeta_L1[23]));
SS_ADDSUB ADDSUB_dbeta_L1_24(.CLK(CLK), .INIT(INIT), .IN({ dbeta_L1_netPar0[24], dbeta_L1_netPar1[24], dbeta_L1_netPar2[24] }), .SIGN({ SIGN_dbeta_L1_netPar0[24], SIGN_dbeta_L1_netPar1[24], SIGN_dbeta_L1_netPar2[24]}), .R_condition(rc[149]), .OUT(dbeta_L1[24]), .SIGN_out(SIGN_dbeta_L1[24]));
defparam ADDSUB_dbeta_L1_0.N = 3;
defparam ADDSUB_dbeta_L1_1.N = 3;
defparam ADDSUB_dbeta_L1_2.N = 3;
defparam ADDSUB_dbeta_L1_3.N = 3;
defparam ADDSUB_dbeta_L1_4.N = 3;
defparam ADDSUB_dbeta_L1_5.N = 3;
defparam ADDSUB_dbeta_L1_6.N = 3;
defparam ADDSUB_dbeta_L1_7.N = 3;
defparam ADDSUB_dbeta_L1_8.N = 3;
defparam ADDSUB_dbeta_L1_9.N = 3;
defparam ADDSUB_dbeta_L1_10.N = 3;
defparam ADDSUB_dbeta_L1_11.N = 3;
defparam ADDSUB_dbeta_L1_12.N = 3;
defparam ADDSUB_dbeta_L1_13.N = 3;
defparam ADDSUB_dbeta_L1_14.N = 3;
defparam ADDSUB_dbeta_L1_15.N = 3;
defparam ADDSUB_dbeta_L1_16.N = 3;
defparam ADDSUB_dbeta_L1_17.N = 3;
defparam ADDSUB_dbeta_L1_18.N = 3;
defparam ADDSUB_dbeta_L1_19.N = 3;
defparam ADDSUB_dbeta_L1_20.N = 3;
defparam ADDSUB_dbeta_L1_21.N = 3;
defparam ADDSUB_dbeta_L1_22.N = 3;
defparam ADDSUB_dbeta_L1_23.N = 3;
defparam ADDSUB_dbeta_L1_24.N = 3;
defparam ADDSUB_dbeta_L1_0.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dbeta_L1_1.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dbeta_L1_2.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dbeta_L1_3.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dbeta_L1_4.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dbeta_L1_5.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dbeta_L1_6.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dbeta_L1_7.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dbeta_L1_8.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dbeta_L1_9.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dbeta_L1_10.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dbeta_L1_11.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dbeta_L1_12.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dbeta_L1_13.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dbeta_L1_14.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dbeta_L1_15.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dbeta_L1_16.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dbeta_L1_17.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dbeta_L1_18.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dbeta_L1_19.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dbeta_L1_20.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dbeta_L1_21.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dbeta_L1_22.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dbeta_L1_23.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dbeta_L1_24.DIFFCOUNTER_SIZE = 3;


SS_ADDSUB ADDSUB_dalpha_L2_0_0(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_0_netPar0[0], dalpha_L2_j_0_netPar1[0], dalpha_L2_j_0_netPar2[0] }), .SIGN({ SIGN_dalpha_L2_j_0_netPar0[0], SIGN_dalpha_L2_j_0_netPar1[0], SIGN_dalpha_L2_j_0_netPar2[0]}), .R_condition(rc[150]), .OUT(dalpha_L2_j_0[0]), .SIGN_out(SIGN_dalpha_L2_j_0[0]));
SS_ADDSUB ADDSUB_dalpha_L2_0_1(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_1_netPar0[0], dalpha_L2_j_1_netPar1[0], dalpha_L2_j_1_netPar2[0] }), .SIGN({ SIGN_dalpha_L2_j_1_netPar0[0], SIGN_dalpha_L2_j_1_netPar1[0], SIGN_dalpha_L2_j_1_netPar2[0]}), .R_condition(rc[151]), .OUT(dalpha_L2_j_1[0]), .SIGN_out(SIGN_dalpha_L2_j_1[0]));
SS_ADDSUB ADDSUB_dalpha_L2_0_2(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_2_netPar0[0], dalpha_L2_j_2_netPar1[0], dalpha_L2_j_2_netPar2[0] }), .SIGN({ SIGN_dalpha_L2_j_2_netPar0[0], SIGN_dalpha_L2_j_2_netPar1[0], SIGN_dalpha_L2_j_2_netPar2[0]}), .R_condition(rc[152]), .OUT(dalpha_L2_j_2[0]), .SIGN_out(SIGN_dalpha_L2_j_2[0]));
SS_ADDSUB ADDSUB_dalpha_L2_0_3(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_3_netPar0[0], dalpha_L2_j_3_netPar1[0], dalpha_L2_j_3_netPar2[0] }), .SIGN({ SIGN_dalpha_L2_j_3_netPar0[0], SIGN_dalpha_L2_j_3_netPar1[0], SIGN_dalpha_L2_j_3_netPar2[0]}), .R_condition(rc[153]), .OUT(dalpha_L2_j_3[0]), .SIGN_out(SIGN_dalpha_L2_j_3[0]));
SS_ADDSUB ADDSUB_dalpha_L2_0_4(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_4_netPar0[0], dalpha_L2_j_4_netPar1[0], dalpha_L2_j_4_netPar2[0] }), .SIGN({ SIGN_dalpha_L2_j_4_netPar0[0], SIGN_dalpha_L2_j_4_netPar1[0], SIGN_dalpha_L2_j_4_netPar2[0]}), .R_condition(rc[154]), .OUT(dalpha_L2_j_4[0]), .SIGN_out(SIGN_dalpha_L2_j_4[0]));
SS_ADDSUB ADDSUB_dalpha_L2_0_5(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_5_netPar0[0], dalpha_L2_j_5_netPar1[0], dalpha_L2_j_5_netPar2[0] }), .SIGN({ SIGN_dalpha_L2_j_5_netPar0[0], SIGN_dalpha_L2_j_5_netPar1[0], SIGN_dalpha_L2_j_5_netPar2[0]}), .R_condition(rc[155]), .OUT(dalpha_L2_j_5[0]), .SIGN_out(SIGN_dalpha_L2_j_5[0]));
SS_ADDSUB ADDSUB_dalpha_L2_0_6(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_6_netPar0[0], dalpha_L2_j_6_netPar1[0], dalpha_L2_j_6_netPar2[0] }), .SIGN({ SIGN_dalpha_L2_j_6_netPar0[0], SIGN_dalpha_L2_j_6_netPar1[0], SIGN_dalpha_L2_j_6_netPar2[0]}), .R_condition(rc[156]), .OUT(dalpha_L2_j_6[0]), .SIGN_out(SIGN_dalpha_L2_j_6[0]));
SS_ADDSUB ADDSUB_dalpha_L2_0_7(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_7_netPar0[0], dalpha_L2_j_7_netPar1[0], dalpha_L2_j_7_netPar2[0] }), .SIGN({ SIGN_dalpha_L2_j_7_netPar0[0], SIGN_dalpha_L2_j_7_netPar1[0], SIGN_dalpha_L2_j_7_netPar2[0]}), .R_condition(rc[157]), .OUT(dalpha_L2_j_7[0]), .SIGN_out(SIGN_dalpha_L2_j_7[0]));
SS_ADDSUB ADDSUB_dalpha_L2_1_0(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_0_netPar0[1], dalpha_L2_j_0_netPar1[1], dalpha_L2_j_0_netPar2[1] }), .SIGN({ SIGN_dalpha_L2_j_0_netPar0[1], SIGN_dalpha_L2_j_0_netPar1[1], SIGN_dalpha_L2_j_0_netPar2[1]}), .R_condition(rc[158]), .OUT(dalpha_L2_j_0[1]), .SIGN_out(SIGN_dalpha_L2_j_0[1]));
SS_ADDSUB ADDSUB_dalpha_L2_1_1(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_1_netPar0[1], dalpha_L2_j_1_netPar1[1], dalpha_L2_j_1_netPar2[1] }), .SIGN({ SIGN_dalpha_L2_j_1_netPar0[1], SIGN_dalpha_L2_j_1_netPar1[1], SIGN_dalpha_L2_j_1_netPar2[1]}), .R_condition(rc[159]), .OUT(dalpha_L2_j_1[1]), .SIGN_out(SIGN_dalpha_L2_j_1[1]));
SS_ADDSUB ADDSUB_dalpha_L2_1_2(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_2_netPar0[1], dalpha_L2_j_2_netPar1[1], dalpha_L2_j_2_netPar2[1] }), .SIGN({ SIGN_dalpha_L2_j_2_netPar0[1], SIGN_dalpha_L2_j_2_netPar1[1], SIGN_dalpha_L2_j_2_netPar2[1]}), .R_condition(rc[160]), .OUT(dalpha_L2_j_2[1]), .SIGN_out(SIGN_dalpha_L2_j_2[1]));
SS_ADDSUB ADDSUB_dalpha_L2_1_3(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_3_netPar0[1], dalpha_L2_j_3_netPar1[1], dalpha_L2_j_3_netPar2[1] }), .SIGN({ SIGN_dalpha_L2_j_3_netPar0[1], SIGN_dalpha_L2_j_3_netPar1[1], SIGN_dalpha_L2_j_3_netPar2[1]}), .R_condition(rc[161]), .OUT(dalpha_L2_j_3[1]), .SIGN_out(SIGN_dalpha_L2_j_3[1]));
SS_ADDSUB ADDSUB_dalpha_L2_1_4(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_4_netPar0[1], dalpha_L2_j_4_netPar1[1], dalpha_L2_j_4_netPar2[1] }), .SIGN({ SIGN_dalpha_L2_j_4_netPar0[1], SIGN_dalpha_L2_j_4_netPar1[1], SIGN_dalpha_L2_j_4_netPar2[1]}), .R_condition(rc[162]), .OUT(dalpha_L2_j_4[1]), .SIGN_out(SIGN_dalpha_L2_j_4[1]));
SS_ADDSUB ADDSUB_dalpha_L2_1_5(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_5_netPar0[1], dalpha_L2_j_5_netPar1[1], dalpha_L2_j_5_netPar2[1] }), .SIGN({ SIGN_dalpha_L2_j_5_netPar0[1], SIGN_dalpha_L2_j_5_netPar1[1], SIGN_dalpha_L2_j_5_netPar2[1]}), .R_condition(rc[163]), .OUT(dalpha_L2_j_5[1]), .SIGN_out(SIGN_dalpha_L2_j_5[1]));
SS_ADDSUB ADDSUB_dalpha_L2_1_6(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_6_netPar0[1], dalpha_L2_j_6_netPar1[1], dalpha_L2_j_6_netPar2[1] }), .SIGN({ SIGN_dalpha_L2_j_6_netPar0[1], SIGN_dalpha_L2_j_6_netPar1[1], SIGN_dalpha_L2_j_6_netPar2[1]}), .R_condition(rc[164]), .OUT(dalpha_L2_j_6[1]), .SIGN_out(SIGN_dalpha_L2_j_6[1]));
SS_ADDSUB ADDSUB_dalpha_L2_1_7(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_7_netPar0[1], dalpha_L2_j_7_netPar1[1], dalpha_L2_j_7_netPar2[1] }), .SIGN({ SIGN_dalpha_L2_j_7_netPar0[1], SIGN_dalpha_L2_j_7_netPar1[1], SIGN_dalpha_L2_j_7_netPar2[1]}), .R_condition(rc[165]), .OUT(dalpha_L2_j_7[1]), .SIGN_out(SIGN_dalpha_L2_j_7[1]));
SS_ADDSUB ADDSUB_dalpha_L2_2_0(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_0_netPar0[2], dalpha_L2_j_0_netPar1[2], dalpha_L2_j_0_netPar2[2] }), .SIGN({ SIGN_dalpha_L2_j_0_netPar0[2], SIGN_dalpha_L2_j_0_netPar1[2], SIGN_dalpha_L2_j_0_netPar2[2]}), .R_condition(rc[166]), .OUT(dalpha_L2_j_0[2]), .SIGN_out(SIGN_dalpha_L2_j_0[2]));
SS_ADDSUB ADDSUB_dalpha_L2_2_1(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_1_netPar0[2], dalpha_L2_j_1_netPar1[2], dalpha_L2_j_1_netPar2[2] }), .SIGN({ SIGN_dalpha_L2_j_1_netPar0[2], SIGN_dalpha_L2_j_1_netPar1[2], SIGN_dalpha_L2_j_1_netPar2[2]}), .R_condition(rc[167]), .OUT(dalpha_L2_j_1[2]), .SIGN_out(SIGN_dalpha_L2_j_1[2]));
SS_ADDSUB ADDSUB_dalpha_L2_2_2(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_2_netPar0[2], dalpha_L2_j_2_netPar1[2], dalpha_L2_j_2_netPar2[2] }), .SIGN({ SIGN_dalpha_L2_j_2_netPar0[2], SIGN_dalpha_L2_j_2_netPar1[2], SIGN_dalpha_L2_j_2_netPar2[2]}), .R_condition(rc[168]), .OUT(dalpha_L2_j_2[2]), .SIGN_out(SIGN_dalpha_L2_j_2[2]));
SS_ADDSUB ADDSUB_dalpha_L2_2_3(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_3_netPar0[2], dalpha_L2_j_3_netPar1[2], dalpha_L2_j_3_netPar2[2] }), .SIGN({ SIGN_dalpha_L2_j_3_netPar0[2], SIGN_dalpha_L2_j_3_netPar1[2], SIGN_dalpha_L2_j_3_netPar2[2]}), .R_condition(rc[169]), .OUT(dalpha_L2_j_3[2]), .SIGN_out(SIGN_dalpha_L2_j_3[2]));
SS_ADDSUB ADDSUB_dalpha_L2_2_4(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_4_netPar0[2], dalpha_L2_j_4_netPar1[2], dalpha_L2_j_4_netPar2[2] }), .SIGN({ SIGN_dalpha_L2_j_4_netPar0[2], SIGN_dalpha_L2_j_4_netPar1[2], SIGN_dalpha_L2_j_4_netPar2[2]}), .R_condition(rc[170]), .OUT(dalpha_L2_j_4[2]), .SIGN_out(SIGN_dalpha_L2_j_4[2]));
SS_ADDSUB ADDSUB_dalpha_L2_2_5(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_5_netPar0[2], dalpha_L2_j_5_netPar1[2], dalpha_L2_j_5_netPar2[2] }), .SIGN({ SIGN_dalpha_L2_j_5_netPar0[2], SIGN_dalpha_L2_j_5_netPar1[2], SIGN_dalpha_L2_j_5_netPar2[2]}), .R_condition(rc[171]), .OUT(dalpha_L2_j_5[2]), .SIGN_out(SIGN_dalpha_L2_j_5[2]));
SS_ADDSUB ADDSUB_dalpha_L2_2_6(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_6_netPar0[2], dalpha_L2_j_6_netPar1[2], dalpha_L2_j_6_netPar2[2] }), .SIGN({ SIGN_dalpha_L2_j_6_netPar0[2], SIGN_dalpha_L2_j_6_netPar1[2], SIGN_dalpha_L2_j_6_netPar2[2]}), .R_condition(rc[172]), .OUT(dalpha_L2_j_6[2]), .SIGN_out(SIGN_dalpha_L2_j_6[2]));
SS_ADDSUB ADDSUB_dalpha_L2_2_7(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_7_netPar0[2], dalpha_L2_j_7_netPar1[2], dalpha_L2_j_7_netPar2[2] }), .SIGN({ SIGN_dalpha_L2_j_7_netPar0[2], SIGN_dalpha_L2_j_7_netPar1[2], SIGN_dalpha_L2_j_7_netPar2[2]}), .R_condition(rc[173]), .OUT(dalpha_L2_j_7[2]), .SIGN_out(SIGN_dalpha_L2_j_7[2]));
SS_ADDSUB ADDSUB_dalpha_L2_3_0(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_0_netPar0[3], dalpha_L2_j_0_netPar1[3], dalpha_L2_j_0_netPar2[3] }), .SIGN({ SIGN_dalpha_L2_j_0_netPar0[3], SIGN_dalpha_L2_j_0_netPar1[3], SIGN_dalpha_L2_j_0_netPar2[3]}), .R_condition(rc[174]), .OUT(dalpha_L2_j_0[3]), .SIGN_out(SIGN_dalpha_L2_j_0[3]));
SS_ADDSUB ADDSUB_dalpha_L2_3_1(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_1_netPar0[3], dalpha_L2_j_1_netPar1[3], dalpha_L2_j_1_netPar2[3] }), .SIGN({ SIGN_dalpha_L2_j_1_netPar0[3], SIGN_dalpha_L2_j_1_netPar1[3], SIGN_dalpha_L2_j_1_netPar2[3]}), .R_condition(rc[175]), .OUT(dalpha_L2_j_1[3]), .SIGN_out(SIGN_dalpha_L2_j_1[3]));
SS_ADDSUB ADDSUB_dalpha_L2_3_2(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_2_netPar0[3], dalpha_L2_j_2_netPar1[3], dalpha_L2_j_2_netPar2[3] }), .SIGN({ SIGN_dalpha_L2_j_2_netPar0[3], SIGN_dalpha_L2_j_2_netPar1[3], SIGN_dalpha_L2_j_2_netPar2[3]}), .R_condition(rc[176]), .OUT(dalpha_L2_j_2[3]), .SIGN_out(SIGN_dalpha_L2_j_2[3]));
SS_ADDSUB ADDSUB_dalpha_L2_3_3(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_3_netPar0[3], dalpha_L2_j_3_netPar1[3], dalpha_L2_j_3_netPar2[3] }), .SIGN({ SIGN_dalpha_L2_j_3_netPar0[3], SIGN_dalpha_L2_j_3_netPar1[3], SIGN_dalpha_L2_j_3_netPar2[3]}), .R_condition(rc[177]), .OUT(dalpha_L2_j_3[3]), .SIGN_out(SIGN_dalpha_L2_j_3[3]));
SS_ADDSUB ADDSUB_dalpha_L2_3_4(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_4_netPar0[3], dalpha_L2_j_4_netPar1[3], dalpha_L2_j_4_netPar2[3] }), .SIGN({ SIGN_dalpha_L2_j_4_netPar0[3], SIGN_dalpha_L2_j_4_netPar1[3], SIGN_dalpha_L2_j_4_netPar2[3]}), .R_condition(rc[178]), .OUT(dalpha_L2_j_4[3]), .SIGN_out(SIGN_dalpha_L2_j_4[3]));
SS_ADDSUB ADDSUB_dalpha_L2_3_5(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_5_netPar0[3], dalpha_L2_j_5_netPar1[3], dalpha_L2_j_5_netPar2[3] }), .SIGN({ SIGN_dalpha_L2_j_5_netPar0[3], SIGN_dalpha_L2_j_5_netPar1[3], SIGN_dalpha_L2_j_5_netPar2[3]}), .R_condition(rc[179]), .OUT(dalpha_L2_j_5[3]), .SIGN_out(SIGN_dalpha_L2_j_5[3]));
SS_ADDSUB ADDSUB_dalpha_L2_3_6(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_6_netPar0[3], dalpha_L2_j_6_netPar1[3], dalpha_L2_j_6_netPar2[3] }), .SIGN({ SIGN_dalpha_L2_j_6_netPar0[3], SIGN_dalpha_L2_j_6_netPar1[3], SIGN_dalpha_L2_j_6_netPar2[3]}), .R_condition(rc[180]), .OUT(dalpha_L2_j_6[3]), .SIGN_out(SIGN_dalpha_L2_j_6[3]));
SS_ADDSUB ADDSUB_dalpha_L2_3_7(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_7_netPar0[3], dalpha_L2_j_7_netPar1[3], dalpha_L2_j_7_netPar2[3] }), .SIGN({ SIGN_dalpha_L2_j_7_netPar0[3], SIGN_dalpha_L2_j_7_netPar1[3], SIGN_dalpha_L2_j_7_netPar2[3]}), .R_condition(rc[181]), .OUT(dalpha_L2_j_7[3]), .SIGN_out(SIGN_dalpha_L2_j_7[3]));
SS_ADDSUB ADDSUB_dalpha_L2_4_0(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_0_netPar0[4], dalpha_L2_j_0_netPar1[4], dalpha_L2_j_0_netPar2[4] }), .SIGN({ SIGN_dalpha_L2_j_0_netPar0[4], SIGN_dalpha_L2_j_0_netPar1[4], SIGN_dalpha_L2_j_0_netPar2[4]}), .R_condition(rc[182]), .OUT(dalpha_L2_j_0[4]), .SIGN_out(SIGN_dalpha_L2_j_0[4]));
SS_ADDSUB ADDSUB_dalpha_L2_4_1(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_1_netPar0[4], dalpha_L2_j_1_netPar1[4], dalpha_L2_j_1_netPar2[4] }), .SIGN({ SIGN_dalpha_L2_j_1_netPar0[4], SIGN_dalpha_L2_j_1_netPar1[4], SIGN_dalpha_L2_j_1_netPar2[4]}), .R_condition(rc[183]), .OUT(dalpha_L2_j_1[4]), .SIGN_out(SIGN_dalpha_L2_j_1[4]));
SS_ADDSUB ADDSUB_dalpha_L2_4_2(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_2_netPar0[4], dalpha_L2_j_2_netPar1[4], dalpha_L2_j_2_netPar2[4] }), .SIGN({ SIGN_dalpha_L2_j_2_netPar0[4], SIGN_dalpha_L2_j_2_netPar1[4], SIGN_dalpha_L2_j_2_netPar2[4]}), .R_condition(rc[184]), .OUT(dalpha_L2_j_2[4]), .SIGN_out(SIGN_dalpha_L2_j_2[4]));
SS_ADDSUB ADDSUB_dalpha_L2_4_3(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_3_netPar0[4], dalpha_L2_j_3_netPar1[4], dalpha_L2_j_3_netPar2[4] }), .SIGN({ SIGN_dalpha_L2_j_3_netPar0[4], SIGN_dalpha_L2_j_3_netPar1[4], SIGN_dalpha_L2_j_3_netPar2[4]}), .R_condition(rc[185]), .OUT(dalpha_L2_j_3[4]), .SIGN_out(SIGN_dalpha_L2_j_3[4]));
SS_ADDSUB ADDSUB_dalpha_L2_4_4(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_4_netPar0[4], dalpha_L2_j_4_netPar1[4], dalpha_L2_j_4_netPar2[4] }), .SIGN({ SIGN_dalpha_L2_j_4_netPar0[4], SIGN_dalpha_L2_j_4_netPar1[4], SIGN_dalpha_L2_j_4_netPar2[4]}), .R_condition(rc[186]), .OUT(dalpha_L2_j_4[4]), .SIGN_out(SIGN_dalpha_L2_j_4[4]));
SS_ADDSUB ADDSUB_dalpha_L2_4_5(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_5_netPar0[4], dalpha_L2_j_5_netPar1[4], dalpha_L2_j_5_netPar2[4] }), .SIGN({ SIGN_dalpha_L2_j_5_netPar0[4], SIGN_dalpha_L2_j_5_netPar1[4], SIGN_dalpha_L2_j_5_netPar2[4]}), .R_condition(rc[187]), .OUT(dalpha_L2_j_5[4]), .SIGN_out(SIGN_dalpha_L2_j_5[4]));
SS_ADDSUB ADDSUB_dalpha_L2_4_6(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_6_netPar0[4], dalpha_L2_j_6_netPar1[4], dalpha_L2_j_6_netPar2[4] }), .SIGN({ SIGN_dalpha_L2_j_6_netPar0[4], SIGN_dalpha_L2_j_6_netPar1[4], SIGN_dalpha_L2_j_6_netPar2[4]}), .R_condition(rc[188]), .OUT(dalpha_L2_j_6[4]), .SIGN_out(SIGN_dalpha_L2_j_6[4]));
SS_ADDSUB ADDSUB_dalpha_L2_4_7(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_7_netPar0[4], dalpha_L2_j_7_netPar1[4], dalpha_L2_j_7_netPar2[4] }), .SIGN({ SIGN_dalpha_L2_j_7_netPar0[4], SIGN_dalpha_L2_j_7_netPar1[4], SIGN_dalpha_L2_j_7_netPar2[4]}), .R_condition(rc[189]), .OUT(dalpha_L2_j_7[4]), .SIGN_out(SIGN_dalpha_L2_j_7[4]));
SS_ADDSUB ADDSUB_dalpha_L2_5_0(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_0_netPar0[5], dalpha_L2_j_0_netPar1[5], dalpha_L2_j_0_netPar2[5] }), .SIGN({ SIGN_dalpha_L2_j_0_netPar0[5], SIGN_dalpha_L2_j_0_netPar1[5], SIGN_dalpha_L2_j_0_netPar2[5]}), .R_condition(rc[190]), .OUT(dalpha_L2_j_0[5]), .SIGN_out(SIGN_dalpha_L2_j_0[5]));
SS_ADDSUB ADDSUB_dalpha_L2_5_1(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_1_netPar0[5], dalpha_L2_j_1_netPar1[5], dalpha_L2_j_1_netPar2[5] }), .SIGN({ SIGN_dalpha_L2_j_1_netPar0[5], SIGN_dalpha_L2_j_1_netPar1[5], SIGN_dalpha_L2_j_1_netPar2[5]}), .R_condition(rc[191]), .OUT(dalpha_L2_j_1[5]), .SIGN_out(SIGN_dalpha_L2_j_1[5]));
SS_ADDSUB ADDSUB_dalpha_L2_5_2(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_2_netPar0[5], dalpha_L2_j_2_netPar1[5], dalpha_L2_j_2_netPar2[5] }), .SIGN({ SIGN_dalpha_L2_j_2_netPar0[5], SIGN_dalpha_L2_j_2_netPar1[5], SIGN_dalpha_L2_j_2_netPar2[5]}), .R_condition(rc[192]), .OUT(dalpha_L2_j_2[5]), .SIGN_out(SIGN_dalpha_L2_j_2[5]));
SS_ADDSUB ADDSUB_dalpha_L2_5_3(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_3_netPar0[5], dalpha_L2_j_3_netPar1[5], dalpha_L2_j_3_netPar2[5] }), .SIGN({ SIGN_dalpha_L2_j_3_netPar0[5], SIGN_dalpha_L2_j_3_netPar1[5], SIGN_dalpha_L2_j_3_netPar2[5]}), .R_condition(rc[193]), .OUT(dalpha_L2_j_3[5]), .SIGN_out(SIGN_dalpha_L2_j_3[5]));
SS_ADDSUB ADDSUB_dalpha_L2_5_4(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_4_netPar0[5], dalpha_L2_j_4_netPar1[5], dalpha_L2_j_4_netPar2[5] }), .SIGN({ SIGN_dalpha_L2_j_4_netPar0[5], SIGN_dalpha_L2_j_4_netPar1[5], SIGN_dalpha_L2_j_4_netPar2[5]}), .R_condition(rc[194]), .OUT(dalpha_L2_j_4[5]), .SIGN_out(SIGN_dalpha_L2_j_4[5]));
SS_ADDSUB ADDSUB_dalpha_L2_5_5(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_5_netPar0[5], dalpha_L2_j_5_netPar1[5], dalpha_L2_j_5_netPar2[5] }), .SIGN({ SIGN_dalpha_L2_j_5_netPar0[5], SIGN_dalpha_L2_j_5_netPar1[5], SIGN_dalpha_L2_j_5_netPar2[5]}), .R_condition(rc[195]), .OUT(dalpha_L2_j_5[5]), .SIGN_out(SIGN_dalpha_L2_j_5[5]));
SS_ADDSUB ADDSUB_dalpha_L2_5_6(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_6_netPar0[5], dalpha_L2_j_6_netPar1[5], dalpha_L2_j_6_netPar2[5] }), .SIGN({ SIGN_dalpha_L2_j_6_netPar0[5], SIGN_dalpha_L2_j_6_netPar1[5], SIGN_dalpha_L2_j_6_netPar2[5]}), .R_condition(rc[196]), .OUT(dalpha_L2_j_6[5]), .SIGN_out(SIGN_dalpha_L2_j_6[5]));
SS_ADDSUB ADDSUB_dalpha_L2_5_7(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_7_netPar0[5], dalpha_L2_j_7_netPar1[5], dalpha_L2_j_7_netPar2[5] }), .SIGN({ SIGN_dalpha_L2_j_7_netPar0[5], SIGN_dalpha_L2_j_7_netPar1[5], SIGN_dalpha_L2_j_7_netPar2[5]}), .R_condition(rc[197]), .OUT(dalpha_L2_j_7[5]), .SIGN_out(SIGN_dalpha_L2_j_7[5]));
SS_ADDSUB ADDSUB_dalpha_L2_6_0(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_0_netPar0[6], dalpha_L2_j_0_netPar1[6], dalpha_L2_j_0_netPar2[6] }), .SIGN({ SIGN_dalpha_L2_j_0_netPar0[6], SIGN_dalpha_L2_j_0_netPar1[6], SIGN_dalpha_L2_j_0_netPar2[6]}), .R_condition(rc[198]), .OUT(dalpha_L2_j_0[6]), .SIGN_out(SIGN_dalpha_L2_j_0[6]));
SS_ADDSUB ADDSUB_dalpha_L2_6_1(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_1_netPar0[6], dalpha_L2_j_1_netPar1[6], dalpha_L2_j_1_netPar2[6] }), .SIGN({ SIGN_dalpha_L2_j_1_netPar0[6], SIGN_dalpha_L2_j_1_netPar1[6], SIGN_dalpha_L2_j_1_netPar2[6]}), .R_condition(rc[199]), .OUT(dalpha_L2_j_1[6]), .SIGN_out(SIGN_dalpha_L2_j_1[6]));
SS_ADDSUB ADDSUB_dalpha_L2_6_2(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_2_netPar0[6], dalpha_L2_j_2_netPar1[6], dalpha_L2_j_2_netPar2[6] }), .SIGN({ SIGN_dalpha_L2_j_2_netPar0[6], SIGN_dalpha_L2_j_2_netPar1[6], SIGN_dalpha_L2_j_2_netPar2[6]}), .R_condition(rc[200]), .OUT(dalpha_L2_j_2[6]), .SIGN_out(SIGN_dalpha_L2_j_2[6]));
SS_ADDSUB ADDSUB_dalpha_L2_6_3(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_3_netPar0[6], dalpha_L2_j_3_netPar1[6], dalpha_L2_j_3_netPar2[6] }), .SIGN({ SIGN_dalpha_L2_j_3_netPar0[6], SIGN_dalpha_L2_j_3_netPar1[6], SIGN_dalpha_L2_j_3_netPar2[6]}), .R_condition(rc[201]), .OUT(dalpha_L2_j_3[6]), .SIGN_out(SIGN_dalpha_L2_j_3[6]));
SS_ADDSUB ADDSUB_dalpha_L2_6_4(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_4_netPar0[6], dalpha_L2_j_4_netPar1[6], dalpha_L2_j_4_netPar2[6] }), .SIGN({ SIGN_dalpha_L2_j_4_netPar0[6], SIGN_dalpha_L2_j_4_netPar1[6], SIGN_dalpha_L2_j_4_netPar2[6]}), .R_condition(rc[202]), .OUT(dalpha_L2_j_4[6]), .SIGN_out(SIGN_dalpha_L2_j_4[6]));
SS_ADDSUB ADDSUB_dalpha_L2_6_5(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_5_netPar0[6], dalpha_L2_j_5_netPar1[6], dalpha_L2_j_5_netPar2[6] }), .SIGN({ SIGN_dalpha_L2_j_5_netPar0[6], SIGN_dalpha_L2_j_5_netPar1[6], SIGN_dalpha_L2_j_5_netPar2[6]}), .R_condition(rc[203]), .OUT(dalpha_L2_j_5[6]), .SIGN_out(SIGN_dalpha_L2_j_5[6]));
SS_ADDSUB ADDSUB_dalpha_L2_6_6(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_6_netPar0[6], dalpha_L2_j_6_netPar1[6], dalpha_L2_j_6_netPar2[6] }), .SIGN({ SIGN_dalpha_L2_j_6_netPar0[6], SIGN_dalpha_L2_j_6_netPar1[6], SIGN_dalpha_L2_j_6_netPar2[6]}), .R_condition(rc[204]), .OUT(dalpha_L2_j_6[6]), .SIGN_out(SIGN_dalpha_L2_j_6[6]));
SS_ADDSUB ADDSUB_dalpha_L2_6_7(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_7_netPar0[6], dalpha_L2_j_7_netPar1[6], dalpha_L2_j_7_netPar2[6] }), .SIGN({ SIGN_dalpha_L2_j_7_netPar0[6], SIGN_dalpha_L2_j_7_netPar1[6], SIGN_dalpha_L2_j_7_netPar2[6]}), .R_condition(rc[205]), .OUT(dalpha_L2_j_7[6]), .SIGN_out(SIGN_dalpha_L2_j_7[6]));
SS_ADDSUB ADDSUB_dalpha_L2_7_0(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_0_netPar0[7], dalpha_L2_j_0_netPar1[7], dalpha_L2_j_0_netPar2[7] }), .SIGN({ SIGN_dalpha_L2_j_0_netPar0[7], SIGN_dalpha_L2_j_0_netPar1[7], SIGN_dalpha_L2_j_0_netPar2[7]}), .R_condition(rc[206]), .OUT(dalpha_L2_j_0[7]), .SIGN_out(SIGN_dalpha_L2_j_0[7]));
SS_ADDSUB ADDSUB_dalpha_L2_7_1(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_1_netPar0[7], dalpha_L2_j_1_netPar1[7], dalpha_L2_j_1_netPar2[7] }), .SIGN({ SIGN_dalpha_L2_j_1_netPar0[7], SIGN_dalpha_L2_j_1_netPar1[7], SIGN_dalpha_L2_j_1_netPar2[7]}), .R_condition(rc[207]), .OUT(dalpha_L2_j_1[7]), .SIGN_out(SIGN_dalpha_L2_j_1[7]));
SS_ADDSUB ADDSUB_dalpha_L2_7_2(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_2_netPar0[7], dalpha_L2_j_2_netPar1[7], dalpha_L2_j_2_netPar2[7] }), .SIGN({ SIGN_dalpha_L2_j_2_netPar0[7], SIGN_dalpha_L2_j_2_netPar1[7], SIGN_dalpha_L2_j_2_netPar2[7]}), .R_condition(rc[208]), .OUT(dalpha_L2_j_2[7]), .SIGN_out(SIGN_dalpha_L2_j_2[7]));
SS_ADDSUB ADDSUB_dalpha_L2_7_3(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_3_netPar0[7], dalpha_L2_j_3_netPar1[7], dalpha_L2_j_3_netPar2[7] }), .SIGN({ SIGN_dalpha_L2_j_3_netPar0[7], SIGN_dalpha_L2_j_3_netPar1[7], SIGN_dalpha_L2_j_3_netPar2[7]}), .R_condition(rc[209]), .OUT(dalpha_L2_j_3[7]), .SIGN_out(SIGN_dalpha_L2_j_3[7]));
SS_ADDSUB ADDSUB_dalpha_L2_7_4(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_4_netPar0[7], dalpha_L2_j_4_netPar1[7], dalpha_L2_j_4_netPar2[7] }), .SIGN({ SIGN_dalpha_L2_j_4_netPar0[7], SIGN_dalpha_L2_j_4_netPar1[7], SIGN_dalpha_L2_j_4_netPar2[7]}), .R_condition(rc[210]), .OUT(dalpha_L2_j_4[7]), .SIGN_out(SIGN_dalpha_L2_j_4[7]));
SS_ADDSUB ADDSUB_dalpha_L2_7_5(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_5_netPar0[7], dalpha_L2_j_5_netPar1[7], dalpha_L2_j_5_netPar2[7] }), .SIGN({ SIGN_dalpha_L2_j_5_netPar0[7], SIGN_dalpha_L2_j_5_netPar1[7], SIGN_dalpha_L2_j_5_netPar2[7]}), .R_condition(rc[211]), .OUT(dalpha_L2_j_5[7]), .SIGN_out(SIGN_dalpha_L2_j_5[7]));
SS_ADDSUB ADDSUB_dalpha_L2_7_6(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_6_netPar0[7], dalpha_L2_j_6_netPar1[7], dalpha_L2_j_6_netPar2[7] }), .SIGN({ SIGN_dalpha_L2_j_6_netPar0[7], SIGN_dalpha_L2_j_6_netPar1[7], SIGN_dalpha_L2_j_6_netPar2[7]}), .R_condition(rc[212]), .OUT(dalpha_L2_j_6[7]), .SIGN_out(SIGN_dalpha_L2_j_6[7]));
SS_ADDSUB ADDSUB_dalpha_L2_7_7(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_7_netPar0[7], dalpha_L2_j_7_netPar1[7], dalpha_L2_j_7_netPar2[7] }), .SIGN({ SIGN_dalpha_L2_j_7_netPar0[7], SIGN_dalpha_L2_j_7_netPar1[7], SIGN_dalpha_L2_j_7_netPar2[7]}), .R_condition(rc[213]), .OUT(dalpha_L2_j_7[7]), .SIGN_out(SIGN_dalpha_L2_j_7[7]));
SS_ADDSUB ADDSUB_dalpha_L2_8_0(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_0_netPar0[8], dalpha_L2_j_0_netPar1[8], dalpha_L2_j_0_netPar2[8] }), .SIGN({ SIGN_dalpha_L2_j_0_netPar0[8], SIGN_dalpha_L2_j_0_netPar1[8], SIGN_dalpha_L2_j_0_netPar2[8]}), .R_condition(rc[214]), .OUT(dalpha_L2_j_0[8]), .SIGN_out(SIGN_dalpha_L2_j_0[8]));
SS_ADDSUB ADDSUB_dalpha_L2_8_1(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_1_netPar0[8], dalpha_L2_j_1_netPar1[8], dalpha_L2_j_1_netPar2[8] }), .SIGN({ SIGN_dalpha_L2_j_1_netPar0[8], SIGN_dalpha_L2_j_1_netPar1[8], SIGN_dalpha_L2_j_1_netPar2[8]}), .R_condition(rc[215]), .OUT(dalpha_L2_j_1[8]), .SIGN_out(SIGN_dalpha_L2_j_1[8]));
SS_ADDSUB ADDSUB_dalpha_L2_8_2(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_2_netPar0[8], dalpha_L2_j_2_netPar1[8], dalpha_L2_j_2_netPar2[8] }), .SIGN({ SIGN_dalpha_L2_j_2_netPar0[8], SIGN_dalpha_L2_j_2_netPar1[8], SIGN_dalpha_L2_j_2_netPar2[8]}), .R_condition(rc[216]), .OUT(dalpha_L2_j_2[8]), .SIGN_out(SIGN_dalpha_L2_j_2[8]));
SS_ADDSUB ADDSUB_dalpha_L2_8_3(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_3_netPar0[8], dalpha_L2_j_3_netPar1[8], dalpha_L2_j_3_netPar2[8] }), .SIGN({ SIGN_dalpha_L2_j_3_netPar0[8], SIGN_dalpha_L2_j_3_netPar1[8], SIGN_dalpha_L2_j_3_netPar2[8]}), .R_condition(rc[217]), .OUT(dalpha_L2_j_3[8]), .SIGN_out(SIGN_dalpha_L2_j_3[8]));
SS_ADDSUB ADDSUB_dalpha_L2_8_4(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_4_netPar0[8], dalpha_L2_j_4_netPar1[8], dalpha_L2_j_4_netPar2[8] }), .SIGN({ SIGN_dalpha_L2_j_4_netPar0[8], SIGN_dalpha_L2_j_4_netPar1[8], SIGN_dalpha_L2_j_4_netPar2[8]}), .R_condition(rc[218]), .OUT(dalpha_L2_j_4[8]), .SIGN_out(SIGN_dalpha_L2_j_4[8]));
SS_ADDSUB ADDSUB_dalpha_L2_8_5(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_5_netPar0[8], dalpha_L2_j_5_netPar1[8], dalpha_L2_j_5_netPar2[8] }), .SIGN({ SIGN_dalpha_L2_j_5_netPar0[8], SIGN_dalpha_L2_j_5_netPar1[8], SIGN_dalpha_L2_j_5_netPar2[8]}), .R_condition(rc[219]), .OUT(dalpha_L2_j_5[8]), .SIGN_out(SIGN_dalpha_L2_j_5[8]));
SS_ADDSUB ADDSUB_dalpha_L2_8_6(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_6_netPar0[8], dalpha_L2_j_6_netPar1[8], dalpha_L2_j_6_netPar2[8] }), .SIGN({ SIGN_dalpha_L2_j_6_netPar0[8], SIGN_dalpha_L2_j_6_netPar1[8], SIGN_dalpha_L2_j_6_netPar2[8]}), .R_condition(rc[220]), .OUT(dalpha_L2_j_6[8]), .SIGN_out(SIGN_dalpha_L2_j_6[8]));
SS_ADDSUB ADDSUB_dalpha_L2_8_7(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_7_netPar0[8], dalpha_L2_j_7_netPar1[8], dalpha_L2_j_7_netPar2[8] }), .SIGN({ SIGN_dalpha_L2_j_7_netPar0[8], SIGN_dalpha_L2_j_7_netPar1[8], SIGN_dalpha_L2_j_7_netPar2[8]}), .R_condition(rc[221]), .OUT(dalpha_L2_j_7[8]), .SIGN_out(SIGN_dalpha_L2_j_7[8]));
SS_ADDSUB ADDSUB_dalpha_L2_9_0(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_0_netPar0[9], dalpha_L2_j_0_netPar1[9], dalpha_L2_j_0_netPar2[9] }), .SIGN({ SIGN_dalpha_L2_j_0_netPar0[9], SIGN_dalpha_L2_j_0_netPar1[9], SIGN_dalpha_L2_j_0_netPar2[9]}), .R_condition(rc[222]), .OUT(dalpha_L2_j_0[9]), .SIGN_out(SIGN_dalpha_L2_j_0[9]));
SS_ADDSUB ADDSUB_dalpha_L2_9_1(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_1_netPar0[9], dalpha_L2_j_1_netPar1[9], dalpha_L2_j_1_netPar2[9] }), .SIGN({ SIGN_dalpha_L2_j_1_netPar0[9], SIGN_dalpha_L2_j_1_netPar1[9], SIGN_dalpha_L2_j_1_netPar2[9]}), .R_condition(rc[223]), .OUT(dalpha_L2_j_1[9]), .SIGN_out(SIGN_dalpha_L2_j_1[9]));
SS_ADDSUB ADDSUB_dalpha_L2_9_2(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_2_netPar0[9], dalpha_L2_j_2_netPar1[9], dalpha_L2_j_2_netPar2[9] }), .SIGN({ SIGN_dalpha_L2_j_2_netPar0[9], SIGN_dalpha_L2_j_2_netPar1[9], SIGN_dalpha_L2_j_2_netPar2[9]}), .R_condition(rc[224]), .OUT(dalpha_L2_j_2[9]), .SIGN_out(SIGN_dalpha_L2_j_2[9]));
SS_ADDSUB ADDSUB_dalpha_L2_9_3(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_3_netPar0[9], dalpha_L2_j_3_netPar1[9], dalpha_L2_j_3_netPar2[9] }), .SIGN({ SIGN_dalpha_L2_j_3_netPar0[9], SIGN_dalpha_L2_j_3_netPar1[9], SIGN_dalpha_L2_j_3_netPar2[9]}), .R_condition(rc[225]), .OUT(dalpha_L2_j_3[9]), .SIGN_out(SIGN_dalpha_L2_j_3[9]));
SS_ADDSUB ADDSUB_dalpha_L2_9_4(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_4_netPar0[9], dalpha_L2_j_4_netPar1[9], dalpha_L2_j_4_netPar2[9] }), .SIGN({ SIGN_dalpha_L2_j_4_netPar0[9], SIGN_dalpha_L2_j_4_netPar1[9], SIGN_dalpha_L2_j_4_netPar2[9]}), .R_condition(rc[226]), .OUT(dalpha_L2_j_4[9]), .SIGN_out(SIGN_dalpha_L2_j_4[9]));
SS_ADDSUB ADDSUB_dalpha_L2_9_5(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_5_netPar0[9], dalpha_L2_j_5_netPar1[9], dalpha_L2_j_5_netPar2[9] }), .SIGN({ SIGN_dalpha_L2_j_5_netPar0[9], SIGN_dalpha_L2_j_5_netPar1[9], SIGN_dalpha_L2_j_5_netPar2[9]}), .R_condition(rc[227]), .OUT(dalpha_L2_j_5[9]), .SIGN_out(SIGN_dalpha_L2_j_5[9]));
SS_ADDSUB ADDSUB_dalpha_L2_9_6(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_6_netPar0[9], dalpha_L2_j_6_netPar1[9], dalpha_L2_j_6_netPar2[9] }), .SIGN({ SIGN_dalpha_L2_j_6_netPar0[9], SIGN_dalpha_L2_j_6_netPar1[9], SIGN_dalpha_L2_j_6_netPar2[9]}), .R_condition(rc[228]), .OUT(dalpha_L2_j_6[9]), .SIGN_out(SIGN_dalpha_L2_j_6[9]));
SS_ADDSUB ADDSUB_dalpha_L2_9_7(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_7_netPar0[9], dalpha_L2_j_7_netPar1[9], dalpha_L2_j_7_netPar2[9] }), .SIGN({ SIGN_dalpha_L2_j_7_netPar0[9], SIGN_dalpha_L2_j_7_netPar1[9], SIGN_dalpha_L2_j_7_netPar2[9]}), .R_condition(rc[229]), .OUT(dalpha_L2_j_7[9]), .SIGN_out(SIGN_dalpha_L2_j_7[9]));
SS_ADDSUB ADDSUB_dalpha_L2_10_0(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_0_netPar0[10], dalpha_L2_j_0_netPar1[10], dalpha_L2_j_0_netPar2[10] }), .SIGN({ SIGN_dalpha_L2_j_0_netPar0[10], SIGN_dalpha_L2_j_0_netPar1[10], SIGN_dalpha_L2_j_0_netPar2[10]}), .R_condition(rc[230]), .OUT(dalpha_L2_j_0[10]), .SIGN_out(SIGN_dalpha_L2_j_0[10]));
SS_ADDSUB ADDSUB_dalpha_L2_10_1(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_1_netPar0[10], dalpha_L2_j_1_netPar1[10], dalpha_L2_j_1_netPar2[10] }), .SIGN({ SIGN_dalpha_L2_j_1_netPar0[10], SIGN_dalpha_L2_j_1_netPar1[10], SIGN_dalpha_L2_j_1_netPar2[10]}), .R_condition(rc[231]), .OUT(dalpha_L2_j_1[10]), .SIGN_out(SIGN_dalpha_L2_j_1[10]));
SS_ADDSUB ADDSUB_dalpha_L2_10_2(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_2_netPar0[10], dalpha_L2_j_2_netPar1[10], dalpha_L2_j_2_netPar2[10] }), .SIGN({ SIGN_dalpha_L2_j_2_netPar0[10], SIGN_dalpha_L2_j_2_netPar1[10], SIGN_dalpha_L2_j_2_netPar2[10]}), .R_condition(rc[232]), .OUT(dalpha_L2_j_2[10]), .SIGN_out(SIGN_dalpha_L2_j_2[10]));
SS_ADDSUB ADDSUB_dalpha_L2_10_3(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_3_netPar0[10], dalpha_L2_j_3_netPar1[10], dalpha_L2_j_3_netPar2[10] }), .SIGN({ SIGN_dalpha_L2_j_3_netPar0[10], SIGN_dalpha_L2_j_3_netPar1[10], SIGN_dalpha_L2_j_3_netPar2[10]}), .R_condition(rc[233]), .OUT(dalpha_L2_j_3[10]), .SIGN_out(SIGN_dalpha_L2_j_3[10]));
SS_ADDSUB ADDSUB_dalpha_L2_10_4(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_4_netPar0[10], dalpha_L2_j_4_netPar1[10], dalpha_L2_j_4_netPar2[10] }), .SIGN({ SIGN_dalpha_L2_j_4_netPar0[10], SIGN_dalpha_L2_j_4_netPar1[10], SIGN_dalpha_L2_j_4_netPar2[10]}), .R_condition(rc[234]), .OUT(dalpha_L2_j_4[10]), .SIGN_out(SIGN_dalpha_L2_j_4[10]));
SS_ADDSUB ADDSUB_dalpha_L2_10_5(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_5_netPar0[10], dalpha_L2_j_5_netPar1[10], dalpha_L2_j_5_netPar2[10] }), .SIGN({ SIGN_dalpha_L2_j_5_netPar0[10], SIGN_dalpha_L2_j_5_netPar1[10], SIGN_dalpha_L2_j_5_netPar2[10]}), .R_condition(rc[235]), .OUT(dalpha_L2_j_5[10]), .SIGN_out(SIGN_dalpha_L2_j_5[10]));
SS_ADDSUB ADDSUB_dalpha_L2_10_6(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_6_netPar0[10], dalpha_L2_j_6_netPar1[10], dalpha_L2_j_6_netPar2[10] }), .SIGN({ SIGN_dalpha_L2_j_6_netPar0[10], SIGN_dalpha_L2_j_6_netPar1[10], SIGN_dalpha_L2_j_6_netPar2[10]}), .R_condition(rc[236]), .OUT(dalpha_L2_j_6[10]), .SIGN_out(SIGN_dalpha_L2_j_6[10]));
SS_ADDSUB ADDSUB_dalpha_L2_10_7(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_7_netPar0[10], dalpha_L2_j_7_netPar1[10], dalpha_L2_j_7_netPar2[10] }), .SIGN({ SIGN_dalpha_L2_j_7_netPar0[10], SIGN_dalpha_L2_j_7_netPar1[10], SIGN_dalpha_L2_j_7_netPar2[10]}), .R_condition(rc[237]), .OUT(dalpha_L2_j_7[10]), .SIGN_out(SIGN_dalpha_L2_j_7[10]));
SS_ADDSUB ADDSUB_dalpha_L2_11_0(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_0_netPar0[11], dalpha_L2_j_0_netPar1[11], dalpha_L2_j_0_netPar2[11] }), .SIGN({ SIGN_dalpha_L2_j_0_netPar0[11], SIGN_dalpha_L2_j_0_netPar1[11], SIGN_dalpha_L2_j_0_netPar2[11]}), .R_condition(rc[238]), .OUT(dalpha_L2_j_0[11]), .SIGN_out(SIGN_dalpha_L2_j_0[11]));
SS_ADDSUB ADDSUB_dalpha_L2_11_1(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_1_netPar0[11], dalpha_L2_j_1_netPar1[11], dalpha_L2_j_1_netPar2[11] }), .SIGN({ SIGN_dalpha_L2_j_1_netPar0[11], SIGN_dalpha_L2_j_1_netPar1[11], SIGN_dalpha_L2_j_1_netPar2[11]}), .R_condition(rc[239]), .OUT(dalpha_L2_j_1[11]), .SIGN_out(SIGN_dalpha_L2_j_1[11]));
SS_ADDSUB ADDSUB_dalpha_L2_11_2(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_2_netPar0[11], dalpha_L2_j_2_netPar1[11], dalpha_L2_j_2_netPar2[11] }), .SIGN({ SIGN_dalpha_L2_j_2_netPar0[11], SIGN_dalpha_L2_j_2_netPar1[11], SIGN_dalpha_L2_j_2_netPar2[11]}), .R_condition(rc[240]), .OUT(dalpha_L2_j_2[11]), .SIGN_out(SIGN_dalpha_L2_j_2[11]));
SS_ADDSUB ADDSUB_dalpha_L2_11_3(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_3_netPar0[11], dalpha_L2_j_3_netPar1[11], dalpha_L2_j_3_netPar2[11] }), .SIGN({ SIGN_dalpha_L2_j_3_netPar0[11], SIGN_dalpha_L2_j_3_netPar1[11], SIGN_dalpha_L2_j_3_netPar2[11]}), .R_condition(rc[241]), .OUT(dalpha_L2_j_3[11]), .SIGN_out(SIGN_dalpha_L2_j_3[11]));
SS_ADDSUB ADDSUB_dalpha_L2_11_4(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_4_netPar0[11], dalpha_L2_j_4_netPar1[11], dalpha_L2_j_4_netPar2[11] }), .SIGN({ SIGN_dalpha_L2_j_4_netPar0[11], SIGN_dalpha_L2_j_4_netPar1[11], SIGN_dalpha_L2_j_4_netPar2[11]}), .R_condition(rc[242]), .OUT(dalpha_L2_j_4[11]), .SIGN_out(SIGN_dalpha_L2_j_4[11]));
SS_ADDSUB ADDSUB_dalpha_L2_11_5(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_5_netPar0[11], dalpha_L2_j_5_netPar1[11], dalpha_L2_j_5_netPar2[11] }), .SIGN({ SIGN_dalpha_L2_j_5_netPar0[11], SIGN_dalpha_L2_j_5_netPar1[11], SIGN_dalpha_L2_j_5_netPar2[11]}), .R_condition(rc[243]), .OUT(dalpha_L2_j_5[11]), .SIGN_out(SIGN_dalpha_L2_j_5[11]));
SS_ADDSUB ADDSUB_dalpha_L2_11_6(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_6_netPar0[11], dalpha_L2_j_6_netPar1[11], dalpha_L2_j_6_netPar2[11] }), .SIGN({ SIGN_dalpha_L2_j_6_netPar0[11], SIGN_dalpha_L2_j_6_netPar1[11], SIGN_dalpha_L2_j_6_netPar2[11]}), .R_condition(rc[244]), .OUT(dalpha_L2_j_6[11]), .SIGN_out(SIGN_dalpha_L2_j_6[11]));
SS_ADDSUB ADDSUB_dalpha_L2_11_7(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_7_netPar0[11], dalpha_L2_j_7_netPar1[11], dalpha_L2_j_7_netPar2[11] }), .SIGN({ SIGN_dalpha_L2_j_7_netPar0[11], SIGN_dalpha_L2_j_7_netPar1[11], SIGN_dalpha_L2_j_7_netPar2[11]}), .R_condition(rc[245]), .OUT(dalpha_L2_j_7[11]), .SIGN_out(SIGN_dalpha_L2_j_7[11]));
SS_ADDSUB ADDSUB_dalpha_L2_12_0(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_0_netPar0[12], dalpha_L2_j_0_netPar1[12], dalpha_L2_j_0_netPar2[12] }), .SIGN({ SIGN_dalpha_L2_j_0_netPar0[12], SIGN_dalpha_L2_j_0_netPar1[12], SIGN_dalpha_L2_j_0_netPar2[12]}), .R_condition(rc[246]), .OUT(dalpha_L2_j_0[12]), .SIGN_out(SIGN_dalpha_L2_j_0[12]));
SS_ADDSUB ADDSUB_dalpha_L2_12_1(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_1_netPar0[12], dalpha_L2_j_1_netPar1[12], dalpha_L2_j_1_netPar2[12] }), .SIGN({ SIGN_dalpha_L2_j_1_netPar0[12], SIGN_dalpha_L2_j_1_netPar1[12], SIGN_dalpha_L2_j_1_netPar2[12]}), .R_condition(rc[247]), .OUT(dalpha_L2_j_1[12]), .SIGN_out(SIGN_dalpha_L2_j_1[12]));
SS_ADDSUB ADDSUB_dalpha_L2_12_2(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_2_netPar0[12], dalpha_L2_j_2_netPar1[12], dalpha_L2_j_2_netPar2[12] }), .SIGN({ SIGN_dalpha_L2_j_2_netPar0[12], SIGN_dalpha_L2_j_2_netPar1[12], SIGN_dalpha_L2_j_2_netPar2[12]}), .R_condition(rc[248]), .OUT(dalpha_L2_j_2[12]), .SIGN_out(SIGN_dalpha_L2_j_2[12]));
SS_ADDSUB ADDSUB_dalpha_L2_12_3(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_3_netPar0[12], dalpha_L2_j_3_netPar1[12], dalpha_L2_j_3_netPar2[12] }), .SIGN({ SIGN_dalpha_L2_j_3_netPar0[12], SIGN_dalpha_L2_j_3_netPar1[12], SIGN_dalpha_L2_j_3_netPar2[12]}), .R_condition(rc[249]), .OUT(dalpha_L2_j_3[12]), .SIGN_out(SIGN_dalpha_L2_j_3[12]));
SS_ADDSUB ADDSUB_dalpha_L2_12_4(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_4_netPar0[12], dalpha_L2_j_4_netPar1[12], dalpha_L2_j_4_netPar2[12] }), .SIGN({ SIGN_dalpha_L2_j_4_netPar0[12], SIGN_dalpha_L2_j_4_netPar1[12], SIGN_dalpha_L2_j_4_netPar2[12]}), .R_condition(rc[250]), .OUT(dalpha_L2_j_4[12]), .SIGN_out(SIGN_dalpha_L2_j_4[12]));
SS_ADDSUB ADDSUB_dalpha_L2_12_5(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_5_netPar0[12], dalpha_L2_j_5_netPar1[12], dalpha_L2_j_5_netPar2[12] }), .SIGN({ SIGN_dalpha_L2_j_5_netPar0[12], SIGN_dalpha_L2_j_5_netPar1[12], SIGN_dalpha_L2_j_5_netPar2[12]}), .R_condition(rc[251]), .OUT(dalpha_L2_j_5[12]), .SIGN_out(SIGN_dalpha_L2_j_5[12]));
SS_ADDSUB ADDSUB_dalpha_L2_12_6(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_6_netPar0[12], dalpha_L2_j_6_netPar1[12], dalpha_L2_j_6_netPar2[12] }), .SIGN({ SIGN_dalpha_L2_j_6_netPar0[12], SIGN_dalpha_L2_j_6_netPar1[12], SIGN_dalpha_L2_j_6_netPar2[12]}), .R_condition(rc[252]), .OUT(dalpha_L2_j_6[12]), .SIGN_out(SIGN_dalpha_L2_j_6[12]));
SS_ADDSUB ADDSUB_dalpha_L2_12_7(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_7_netPar0[12], dalpha_L2_j_7_netPar1[12], dalpha_L2_j_7_netPar2[12] }), .SIGN({ SIGN_dalpha_L2_j_7_netPar0[12], SIGN_dalpha_L2_j_7_netPar1[12], SIGN_dalpha_L2_j_7_netPar2[12]}), .R_condition(rc[253]), .OUT(dalpha_L2_j_7[12]), .SIGN_out(SIGN_dalpha_L2_j_7[12]));
SS_ADDSUB ADDSUB_dalpha_L2_13_0(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_0_netPar0[13], dalpha_L2_j_0_netPar1[13], dalpha_L2_j_0_netPar2[13] }), .SIGN({ SIGN_dalpha_L2_j_0_netPar0[13], SIGN_dalpha_L2_j_0_netPar1[13], SIGN_dalpha_L2_j_0_netPar2[13]}), .R_condition(rc[254]), .OUT(dalpha_L2_j_0[13]), .SIGN_out(SIGN_dalpha_L2_j_0[13]));
SS_ADDSUB ADDSUB_dalpha_L2_13_1(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_1_netPar0[13], dalpha_L2_j_1_netPar1[13], dalpha_L2_j_1_netPar2[13] }), .SIGN({ SIGN_dalpha_L2_j_1_netPar0[13], SIGN_dalpha_L2_j_1_netPar1[13], SIGN_dalpha_L2_j_1_netPar2[13]}), .R_condition(rc[255]), .OUT(dalpha_L2_j_1[13]), .SIGN_out(SIGN_dalpha_L2_j_1[13]));
SS_ADDSUB ADDSUB_dalpha_L2_13_2(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_2_netPar0[13], dalpha_L2_j_2_netPar1[13], dalpha_L2_j_2_netPar2[13] }), .SIGN({ SIGN_dalpha_L2_j_2_netPar0[13], SIGN_dalpha_L2_j_2_netPar1[13], SIGN_dalpha_L2_j_2_netPar2[13]}), .R_condition(rc[256]), .OUT(dalpha_L2_j_2[13]), .SIGN_out(SIGN_dalpha_L2_j_2[13]));
SS_ADDSUB ADDSUB_dalpha_L2_13_3(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_3_netPar0[13], dalpha_L2_j_3_netPar1[13], dalpha_L2_j_3_netPar2[13] }), .SIGN({ SIGN_dalpha_L2_j_3_netPar0[13], SIGN_dalpha_L2_j_3_netPar1[13], SIGN_dalpha_L2_j_3_netPar2[13]}), .R_condition(rc[257]), .OUT(dalpha_L2_j_3[13]), .SIGN_out(SIGN_dalpha_L2_j_3[13]));
SS_ADDSUB ADDSUB_dalpha_L2_13_4(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_4_netPar0[13], dalpha_L2_j_4_netPar1[13], dalpha_L2_j_4_netPar2[13] }), .SIGN({ SIGN_dalpha_L2_j_4_netPar0[13], SIGN_dalpha_L2_j_4_netPar1[13], SIGN_dalpha_L2_j_4_netPar2[13]}), .R_condition(rc[258]), .OUT(dalpha_L2_j_4[13]), .SIGN_out(SIGN_dalpha_L2_j_4[13]));
SS_ADDSUB ADDSUB_dalpha_L2_13_5(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_5_netPar0[13], dalpha_L2_j_5_netPar1[13], dalpha_L2_j_5_netPar2[13] }), .SIGN({ SIGN_dalpha_L2_j_5_netPar0[13], SIGN_dalpha_L2_j_5_netPar1[13], SIGN_dalpha_L2_j_5_netPar2[13]}), .R_condition(rc[259]), .OUT(dalpha_L2_j_5[13]), .SIGN_out(SIGN_dalpha_L2_j_5[13]));
SS_ADDSUB ADDSUB_dalpha_L2_13_6(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_6_netPar0[13], dalpha_L2_j_6_netPar1[13], dalpha_L2_j_6_netPar2[13] }), .SIGN({ SIGN_dalpha_L2_j_6_netPar0[13], SIGN_dalpha_L2_j_6_netPar1[13], SIGN_dalpha_L2_j_6_netPar2[13]}), .R_condition(rc[260]), .OUT(dalpha_L2_j_6[13]), .SIGN_out(SIGN_dalpha_L2_j_6[13]));
SS_ADDSUB ADDSUB_dalpha_L2_13_7(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_7_netPar0[13], dalpha_L2_j_7_netPar1[13], dalpha_L2_j_7_netPar2[13] }), .SIGN({ SIGN_dalpha_L2_j_7_netPar0[13], SIGN_dalpha_L2_j_7_netPar1[13], SIGN_dalpha_L2_j_7_netPar2[13]}), .R_condition(rc[261]), .OUT(dalpha_L2_j_7[13]), .SIGN_out(SIGN_dalpha_L2_j_7[13]));
SS_ADDSUB ADDSUB_dalpha_L2_14_0(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_0_netPar0[14], dalpha_L2_j_0_netPar1[14], dalpha_L2_j_0_netPar2[14] }), .SIGN({ SIGN_dalpha_L2_j_0_netPar0[14], SIGN_dalpha_L2_j_0_netPar1[14], SIGN_dalpha_L2_j_0_netPar2[14]}), .R_condition(rc[262]), .OUT(dalpha_L2_j_0[14]), .SIGN_out(SIGN_dalpha_L2_j_0[14]));
SS_ADDSUB ADDSUB_dalpha_L2_14_1(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_1_netPar0[14], dalpha_L2_j_1_netPar1[14], dalpha_L2_j_1_netPar2[14] }), .SIGN({ SIGN_dalpha_L2_j_1_netPar0[14], SIGN_dalpha_L2_j_1_netPar1[14], SIGN_dalpha_L2_j_1_netPar2[14]}), .R_condition(rc[263]), .OUT(dalpha_L2_j_1[14]), .SIGN_out(SIGN_dalpha_L2_j_1[14]));
SS_ADDSUB ADDSUB_dalpha_L2_14_2(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_2_netPar0[14], dalpha_L2_j_2_netPar1[14], dalpha_L2_j_2_netPar2[14] }), .SIGN({ SIGN_dalpha_L2_j_2_netPar0[14], SIGN_dalpha_L2_j_2_netPar1[14], SIGN_dalpha_L2_j_2_netPar2[14]}), .R_condition(rc[264]), .OUT(dalpha_L2_j_2[14]), .SIGN_out(SIGN_dalpha_L2_j_2[14]));
SS_ADDSUB ADDSUB_dalpha_L2_14_3(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_3_netPar0[14], dalpha_L2_j_3_netPar1[14], dalpha_L2_j_3_netPar2[14] }), .SIGN({ SIGN_dalpha_L2_j_3_netPar0[14], SIGN_dalpha_L2_j_3_netPar1[14], SIGN_dalpha_L2_j_3_netPar2[14]}), .R_condition(rc[265]), .OUT(dalpha_L2_j_3[14]), .SIGN_out(SIGN_dalpha_L2_j_3[14]));
SS_ADDSUB ADDSUB_dalpha_L2_14_4(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_4_netPar0[14], dalpha_L2_j_4_netPar1[14], dalpha_L2_j_4_netPar2[14] }), .SIGN({ SIGN_dalpha_L2_j_4_netPar0[14], SIGN_dalpha_L2_j_4_netPar1[14], SIGN_dalpha_L2_j_4_netPar2[14]}), .R_condition(rc[266]), .OUT(dalpha_L2_j_4[14]), .SIGN_out(SIGN_dalpha_L2_j_4[14]));
SS_ADDSUB ADDSUB_dalpha_L2_14_5(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_5_netPar0[14], dalpha_L2_j_5_netPar1[14], dalpha_L2_j_5_netPar2[14] }), .SIGN({ SIGN_dalpha_L2_j_5_netPar0[14], SIGN_dalpha_L2_j_5_netPar1[14], SIGN_dalpha_L2_j_5_netPar2[14]}), .R_condition(rc[267]), .OUT(dalpha_L2_j_5[14]), .SIGN_out(SIGN_dalpha_L2_j_5[14]));
SS_ADDSUB ADDSUB_dalpha_L2_14_6(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_6_netPar0[14], dalpha_L2_j_6_netPar1[14], dalpha_L2_j_6_netPar2[14] }), .SIGN({ SIGN_dalpha_L2_j_6_netPar0[14], SIGN_dalpha_L2_j_6_netPar1[14], SIGN_dalpha_L2_j_6_netPar2[14]}), .R_condition(rc[268]), .OUT(dalpha_L2_j_6[14]), .SIGN_out(SIGN_dalpha_L2_j_6[14]));
SS_ADDSUB ADDSUB_dalpha_L2_14_7(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_7_netPar0[14], dalpha_L2_j_7_netPar1[14], dalpha_L2_j_7_netPar2[14] }), .SIGN({ SIGN_dalpha_L2_j_7_netPar0[14], SIGN_dalpha_L2_j_7_netPar1[14], SIGN_dalpha_L2_j_7_netPar2[14]}), .R_condition(rc[269]), .OUT(dalpha_L2_j_7[14]), .SIGN_out(SIGN_dalpha_L2_j_7[14]));
SS_ADDSUB ADDSUB_dalpha_L2_15_0(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_0_netPar0[15], dalpha_L2_j_0_netPar1[15], dalpha_L2_j_0_netPar2[15] }), .SIGN({ SIGN_dalpha_L2_j_0_netPar0[15], SIGN_dalpha_L2_j_0_netPar1[15], SIGN_dalpha_L2_j_0_netPar2[15]}), .R_condition(rc[270]), .OUT(dalpha_L2_j_0[15]), .SIGN_out(SIGN_dalpha_L2_j_0[15]));
SS_ADDSUB ADDSUB_dalpha_L2_15_1(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_1_netPar0[15], dalpha_L2_j_1_netPar1[15], dalpha_L2_j_1_netPar2[15] }), .SIGN({ SIGN_dalpha_L2_j_1_netPar0[15], SIGN_dalpha_L2_j_1_netPar1[15], SIGN_dalpha_L2_j_1_netPar2[15]}), .R_condition(rc[271]), .OUT(dalpha_L2_j_1[15]), .SIGN_out(SIGN_dalpha_L2_j_1[15]));
SS_ADDSUB ADDSUB_dalpha_L2_15_2(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_2_netPar0[15], dalpha_L2_j_2_netPar1[15], dalpha_L2_j_2_netPar2[15] }), .SIGN({ SIGN_dalpha_L2_j_2_netPar0[15], SIGN_dalpha_L2_j_2_netPar1[15], SIGN_dalpha_L2_j_2_netPar2[15]}), .R_condition(rc[272]), .OUT(dalpha_L2_j_2[15]), .SIGN_out(SIGN_dalpha_L2_j_2[15]));
SS_ADDSUB ADDSUB_dalpha_L2_15_3(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_3_netPar0[15], dalpha_L2_j_3_netPar1[15], dalpha_L2_j_3_netPar2[15] }), .SIGN({ SIGN_dalpha_L2_j_3_netPar0[15], SIGN_dalpha_L2_j_3_netPar1[15], SIGN_dalpha_L2_j_3_netPar2[15]}), .R_condition(rc[273]), .OUT(dalpha_L2_j_3[15]), .SIGN_out(SIGN_dalpha_L2_j_3[15]));
SS_ADDSUB ADDSUB_dalpha_L2_15_4(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_4_netPar0[15], dalpha_L2_j_4_netPar1[15], dalpha_L2_j_4_netPar2[15] }), .SIGN({ SIGN_dalpha_L2_j_4_netPar0[15], SIGN_dalpha_L2_j_4_netPar1[15], SIGN_dalpha_L2_j_4_netPar2[15]}), .R_condition(rc[274]), .OUT(dalpha_L2_j_4[15]), .SIGN_out(SIGN_dalpha_L2_j_4[15]));
SS_ADDSUB ADDSUB_dalpha_L2_15_5(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_5_netPar0[15], dalpha_L2_j_5_netPar1[15], dalpha_L2_j_5_netPar2[15] }), .SIGN({ SIGN_dalpha_L2_j_5_netPar0[15], SIGN_dalpha_L2_j_5_netPar1[15], SIGN_dalpha_L2_j_5_netPar2[15]}), .R_condition(rc[275]), .OUT(dalpha_L2_j_5[15]), .SIGN_out(SIGN_dalpha_L2_j_5[15]));
SS_ADDSUB ADDSUB_dalpha_L2_15_6(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_6_netPar0[15], dalpha_L2_j_6_netPar1[15], dalpha_L2_j_6_netPar2[15] }), .SIGN({ SIGN_dalpha_L2_j_6_netPar0[15], SIGN_dalpha_L2_j_6_netPar1[15], SIGN_dalpha_L2_j_6_netPar2[15]}), .R_condition(rc[276]), .OUT(dalpha_L2_j_6[15]), .SIGN_out(SIGN_dalpha_L2_j_6[15]));
SS_ADDSUB ADDSUB_dalpha_L2_15_7(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_7_netPar0[15], dalpha_L2_j_7_netPar1[15], dalpha_L2_j_7_netPar2[15] }), .SIGN({ SIGN_dalpha_L2_j_7_netPar0[15], SIGN_dalpha_L2_j_7_netPar1[15], SIGN_dalpha_L2_j_7_netPar2[15]}), .R_condition(rc[277]), .OUT(dalpha_L2_j_7[15]), .SIGN_out(SIGN_dalpha_L2_j_7[15]));
SS_ADDSUB ADDSUB_dalpha_L2_16_0(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_0_netPar0[16], dalpha_L2_j_0_netPar1[16], dalpha_L2_j_0_netPar2[16] }), .SIGN({ SIGN_dalpha_L2_j_0_netPar0[16], SIGN_dalpha_L2_j_0_netPar1[16], SIGN_dalpha_L2_j_0_netPar2[16]}), .R_condition(rc[278]), .OUT(dalpha_L2_j_0[16]), .SIGN_out(SIGN_dalpha_L2_j_0[16]));
SS_ADDSUB ADDSUB_dalpha_L2_16_1(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_1_netPar0[16], dalpha_L2_j_1_netPar1[16], dalpha_L2_j_1_netPar2[16] }), .SIGN({ SIGN_dalpha_L2_j_1_netPar0[16], SIGN_dalpha_L2_j_1_netPar1[16], SIGN_dalpha_L2_j_1_netPar2[16]}), .R_condition(rc[279]), .OUT(dalpha_L2_j_1[16]), .SIGN_out(SIGN_dalpha_L2_j_1[16]));
SS_ADDSUB ADDSUB_dalpha_L2_16_2(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_2_netPar0[16], dalpha_L2_j_2_netPar1[16], dalpha_L2_j_2_netPar2[16] }), .SIGN({ SIGN_dalpha_L2_j_2_netPar0[16], SIGN_dalpha_L2_j_2_netPar1[16], SIGN_dalpha_L2_j_2_netPar2[16]}), .R_condition(rc[280]), .OUT(dalpha_L2_j_2[16]), .SIGN_out(SIGN_dalpha_L2_j_2[16]));
SS_ADDSUB ADDSUB_dalpha_L2_16_3(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_3_netPar0[16], dalpha_L2_j_3_netPar1[16], dalpha_L2_j_3_netPar2[16] }), .SIGN({ SIGN_dalpha_L2_j_3_netPar0[16], SIGN_dalpha_L2_j_3_netPar1[16], SIGN_dalpha_L2_j_3_netPar2[16]}), .R_condition(rc[281]), .OUT(dalpha_L2_j_3[16]), .SIGN_out(SIGN_dalpha_L2_j_3[16]));
SS_ADDSUB ADDSUB_dalpha_L2_16_4(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_4_netPar0[16], dalpha_L2_j_4_netPar1[16], dalpha_L2_j_4_netPar2[16] }), .SIGN({ SIGN_dalpha_L2_j_4_netPar0[16], SIGN_dalpha_L2_j_4_netPar1[16], SIGN_dalpha_L2_j_4_netPar2[16]}), .R_condition(rc[282]), .OUT(dalpha_L2_j_4[16]), .SIGN_out(SIGN_dalpha_L2_j_4[16]));
SS_ADDSUB ADDSUB_dalpha_L2_16_5(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_5_netPar0[16], dalpha_L2_j_5_netPar1[16], dalpha_L2_j_5_netPar2[16] }), .SIGN({ SIGN_dalpha_L2_j_5_netPar0[16], SIGN_dalpha_L2_j_5_netPar1[16], SIGN_dalpha_L2_j_5_netPar2[16]}), .R_condition(rc[283]), .OUT(dalpha_L2_j_5[16]), .SIGN_out(SIGN_dalpha_L2_j_5[16]));
SS_ADDSUB ADDSUB_dalpha_L2_16_6(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_6_netPar0[16], dalpha_L2_j_6_netPar1[16], dalpha_L2_j_6_netPar2[16] }), .SIGN({ SIGN_dalpha_L2_j_6_netPar0[16], SIGN_dalpha_L2_j_6_netPar1[16], SIGN_dalpha_L2_j_6_netPar2[16]}), .R_condition(rc[284]), .OUT(dalpha_L2_j_6[16]), .SIGN_out(SIGN_dalpha_L2_j_6[16]));
SS_ADDSUB ADDSUB_dalpha_L2_16_7(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_7_netPar0[16], dalpha_L2_j_7_netPar1[16], dalpha_L2_j_7_netPar2[16] }), .SIGN({ SIGN_dalpha_L2_j_7_netPar0[16], SIGN_dalpha_L2_j_7_netPar1[16], SIGN_dalpha_L2_j_7_netPar2[16]}), .R_condition(rc[285]), .OUT(dalpha_L2_j_7[16]), .SIGN_out(SIGN_dalpha_L2_j_7[16]));
SS_ADDSUB ADDSUB_dalpha_L2_17_0(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_0_netPar0[17], dalpha_L2_j_0_netPar1[17], dalpha_L2_j_0_netPar2[17] }), .SIGN({ SIGN_dalpha_L2_j_0_netPar0[17], SIGN_dalpha_L2_j_0_netPar1[17], SIGN_dalpha_L2_j_0_netPar2[17]}), .R_condition(rc[286]), .OUT(dalpha_L2_j_0[17]), .SIGN_out(SIGN_dalpha_L2_j_0[17]));
SS_ADDSUB ADDSUB_dalpha_L2_17_1(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_1_netPar0[17], dalpha_L2_j_1_netPar1[17], dalpha_L2_j_1_netPar2[17] }), .SIGN({ SIGN_dalpha_L2_j_1_netPar0[17], SIGN_dalpha_L2_j_1_netPar1[17], SIGN_dalpha_L2_j_1_netPar2[17]}), .R_condition(rc[287]), .OUT(dalpha_L2_j_1[17]), .SIGN_out(SIGN_dalpha_L2_j_1[17]));
SS_ADDSUB ADDSUB_dalpha_L2_17_2(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_2_netPar0[17], dalpha_L2_j_2_netPar1[17], dalpha_L2_j_2_netPar2[17] }), .SIGN({ SIGN_dalpha_L2_j_2_netPar0[17], SIGN_dalpha_L2_j_2_netPar1[17], SIGN_dalpha_L2_j_2_netPar2[17]}), .R_condition(rc[288]), .OUT(dalpha_L2_j_2[17]), .SIGN_out(SIGN_dalpha_L2_j_2[17]));
SS_ADDSUB ADDSUB_dalpha_L2_17_3(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_3_netPar0[17], dalpha_L2_j_3_netPar1[17], dalpha_L2_j_3_netPar2[17] }), .SIGN({ SIGN_dalpha_L2_j_3_netPar0[17], SIGN_dalpha_L2_j_3_netPar1[17], SIGN_dalpha_L2_j_3_netPar2[17]}), .R_condition(rc[289]), .OUT(dalpha_L2_j_3[17]), .SIGN_out(SIGN_dalpha_L2_j_3[17]));
SS_ADDSUB ADDSUB_dalpha_L2_17_4(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_4_netPar0[17], dalpha_L2_j_4_netPar1[17], dalpha_L2_j_4_netPar2[17] }), .SIGN({ SIGN_dalpha_L2_j_4_netPar0[17], SIGN_dalpha_L2_j_4_netPar1[17], SIGN_dalpha_L2_j_4_netPar2[17]}), .R_condition(rc[290]), .OUT(dalpha_L2_j_4[17]), .SIGN_out(SIGN_dalpha_L2_j_4[17]));
SS_ADDSUB ADDSUB_dalpha_L2_17_5(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_5_netPar0[17], dalpha_L2_j_5_netPar1[17], dalpha_L2_j_5_netPar2[17] }), .SIGN({ SIGN_dalpha_L2_j_5_netPar0[17], SIGN_dalpha_L2_j_5_netPar1[17], SIGN_dalpha_L2_j_5_netPar2[17]}), .R_condition(rc[291]), .OUT(dalpha_L2_j_5[17]), .SIGN_out(SIGN_dalpha_L2_j_5[17]));
SS_ADDSUB ADDSUB_dalpha_L2_17_6(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_6_netPar0[17], dalpha_L2_j_6_netPar1[17], dalpha_L2_j_6_netPar2[17] }), .SIGN({ SIGN_dalpha_L2_j_6_netPar0[17], SIGN_dalpha_L2_j_6_netPar1[17], SIGN_dalpha_L2_j_6_netPar2[17]}), .R_condition(rc[292]), .OUT(dalpha_L2_j_6[17]), .SIGN_out(SIGN_dalpha_L2_j_6[17]));
SS_ADDSUB ADDSUB_dalpha_L2_17_7(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_7_netPar0[17], dalpha_L2_j_7_netPar1[17], dalpha_L2_j_7_netPar2[17] }), .SIGN({ SIGN_dalpha_L2_j_7_netPar0[17], SIGN_dalpha_L2_j_7_netPar1[17], SIGN_dalpha_L2_j_7_netPar2[17]}), .R_condition(rc[293]), .OUT(dalpha_L2_j_7[17]), .SIGN_out(SIGN_dalpha_L2_j_7[17]));
SS_ADDSUB ADDSUB_dalpha_L2_18_0(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_0_netPar0[18], dalpha_L2_j_0_netPar1[18], dalpha_L2_j_0_netPar2[18] }), .SIGN({ SIGN_dalpha_L2_j_0_netPar0[18], SIGN_dalpha_L2_j_0_netPar1[18], SIGN_dalpha_L2_j_0_netPar2[18]}), .R_condition(rc[294]), .OUT(dalpha_L2_j_0[18]), .SIGN_out(SIGN_dalpha_L2_j_0[18]));
SS_ADDSUB ADDSUB_dalpha_L2_18_1(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_1_netPar0[18], dalpha_L2_j_1_netPar1[18], dalpha_L2_j_1_netPar2[18] }), .SIGN({ SIGN_dalpha_L2_j_1_netPar0[18], SIGN_dalpha_L2_j_1_netPar1[18], SIGN_dalpha_L2_j_1_netPar2[18]}), .R_condition(rc[295]), .OUT(dalpha_L2_j_1[18]), .SIGN_out(SIGN_dalpha_L2_j_1[18]));
SS_ADDSUB ADDSUB_dalpha_L2_18_2(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_2_netPar0[18], dalpha_L2_j_2_netPar1[18], dalpha_L2_j_2_netPar2[18] }), .SIGN({ SIGN_dalpha_L2_j_2_netPar0[18], SIGN_dalpha_L2_j_2_netPar1[18], SIGN_dalpha_L2_j_2_netPar2[18]}), .R_condition(rc[296]), .OUT(dalpha_L2_j_2[18]), .SIGN_out(SIGN_dalpha_L2_j_2[18]));
SS_ADDSUB ADDSUB_dalpha_L2_18_3(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_3_netPar0[18], dalpha_L2_j_3_netPar1[18], dalpha_L2_j_3_netPar2[18] }), .SIGN({ SIGN_dalpha_L2_j_3_netPar0[18], SIGN_dalpha_L2_j_3_netPar1[18], SIGN_dalpha_L2_j_3_netPar2[18]}), .R_condition(rc[297]), .OUT(dalpha_L2_j_3[18]), .SIGN_out(SIGN_dalpha_L2_j_3[18]));
SS_ADDSUB ADDSUB_dalpha_L2_18_4(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_4_netPar0[18], dalpha_L2_j_4_netPar1[18], dalpha_L2_j_4_netPar2[18] }), .SIGN({ SIGN_dalpha_L2_j_4_netPar0[18], SIGN_dalpha_L2_j_4_netPar1[18], SIGN_dalpha_L2_j_4_netPar2[18]}), .R_condition(rc[298]), .OUT(dalpha_L2_j_4[18]), .SIGN_out(SIGN_dalpha_L2_j_4[18]));
SS_ADDSUB ADDSUB_dalpha_L2_18_5(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_5_netPar0[18], dalpha_L2_j_5_netPar1[18], dalpha_L2_j_5_netPar2[18] }), .SIGN({ SIGN_dalpha_L2_j_5_netPar0[18], SIGN_dalpha_L2_j_5_netPar1[18], SIGN_dalpha_L2_j_5_netPar2[18]}), .R_condition(rc[299]), .OUT(dalpha_L2_j_5[18]), .SIGN_out(SIGN_dalpha_L2_j_5[18]));
SS_ADDSUB ADDSUB_dalpha_L2_18_6(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_6_netPar0[18], dalpha_L2_j_6_netPar1[18], dalpha_L2_j_6_netPar2[18] }), .SIGN({ SIGN_dalpha_L2_j_6_netPar0[18], SIGN_dalpha_L2_j_6_netPar1[18], SIGN_dalpha_L2_j_6_netPar2[18]}), .R_condition(rc[300]), .OUT(dalpha_L2_j_6[18]), .SIGN_out(SIGN_dalpha_L2_j_6[18]));
SS_ADDSUB ADDSUB_dalpha_L2_18_7(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_7_netPar0[18], dalpha_L2_j_7_netPar1[18], dalpha_L2_j_7_netPar2[18] }), .SIGN({ SIGN_dalpha_L2_j_7_netPar0[18], SIGN_dalpha_L2_j_7_netPar1[18], SIGN_dalpha_L2_j_7_netPar2[18]}), .R_condition(rc[301]), .OUT(dalpha_L2_j_7[18]), .SIGN_out(SIGN_dalpha_L2_j_7[18]));
SS_ADDSUB ADDSUB_dalpha_L2_19_0(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_0_netPar0[19], dalpha_L2_j_0_netPar1[19], dalpha_L2_j_0_netPar2[19] }), .SIGN({ SIGN_dalpha_L2_j_0_netPar0[19], SIGN_dalpha_L2_j_0_netPar1[19], SIGN_dalpha_L2_j_0_netPar2[19]}), .R_condition(rc[302]), .OUT(dalpha_L2_j_0[19]), .SIGN_out(SIGN_dalpha_L2_j_0[19]));
SS_ADDSUB ADDSUB_dalpha_L2_19_1(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_1_netPar0[19], dalpha_L2_j_1_netPar1[19], dalpha_L2_j_1_netPar2[19] }), .SIGN({ SIGN_dalpha_L2_j_1_netPar0[19], SIGN_dalpha_L2_j_1_netPar1[19], SIGN_dalpha_L2_j_1_netPar2[19]}), .R_condition(rc[303]), .OUT(dalpha_L2_j_1[19]), .SIGN_out(SIGN_dalpha_L2_j_1[19]));
SS_ADDSUB ADDSUB_dalpha_L2_19_2(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_2_netPar0[19], dalpha_L2_j_2_netPar1[19], dalpha_L2_j_2_netPar2[19] }), .SIGN({ SIGN_dalpha_L2_j_2_netPar0[19], SIGN_dalpha_L2_j_2_netPar1[19], SIGN_dalpha_L2_j_2_netPar2[19]}), .R_condition(rc[304]), .OUT(dalpha_L2_j_2[19]), .SIGN_out(SIGN_dalpha_L2_j_2[19]));
SS_ADDSUB ADDSUB_dalpha_L2_19_3(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_3_netPar0[19], dalpha_L2_j_3_netPar1[19], dalpha_L2_j_3_netPar2[19] }), .SIGN({ SIGN_dalpha_L2_j_3_netPar0[19], SIGN_dalpha_L2_j_3_netPar1[19], SIGN_dalpha_L2_j_3_netPar2[19]}), .R_condition(rc[305]), .OUT(dalpha_L2_j_3[19]), .SIGN_out(SIGN_dalpha_L2_j_3[19]));
SS_ADDSUB ADDSUB_dalpha_L2_19_4(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_4_netPar0[19], dalpha_L2_j_4_netPar1[19], dalpha_L2_j_4_netPar2[19] }), .SIGN({ SIGN_dalpha_L2_j_4_netPar0[19], SIGN_dalpha_L2_j_4_netPar1[19], SIGN_dalpha_L2_j_4_netPar2[19]}), .R_condition(rc[306]), .OUT(dalpha_L2_j_4[19]), .SIGN_out(SIGN_dalpha_L2_j_4[19]));
SS_ADDSUB ADDSUB_dalpha_L2_19_5(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_5_netPar0[19], dalpha_L2_j_5_netPar1[19], dalpha_L2_j_5_netPar2[19] }), .SIGN({ SIGN_dalpha_L2_j_5_netPar0[19], SIGN_dalpha_L2_j_5_netPar1[19], SIGN_dalpha_L2_j_5_netPar2[19]}), .R_condition(rc[307]), .OUT(dalpha_L2_j_5[19]), .SIGN_out(SIGN_dalpha_L2_j_5[19]));
SS_ADDSUB ADDSUB_dalpha_L2_19_6(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_6_netPar0[19], dalpha_L2_j_6_netPar1[19], dalpha_L2_j_6_netPar2[19] }), .SIGN({ SIGN_dalpha_L2_j_6_netPar0[19], SIGN_dalpha_L2_j_6_netPar1[19], SIGN_dalpha_L2_j_6_netPar2[19]}), .R_condition(rc[308]), .OUT(dalpha_L2_j_6[19]), .SIGN_out(SIGN_dalpha_L2_j_6[19]));
SS_ADDSUB ADDSUB_dalpha_L2_19_7(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_7_netPar0[19], dalpha_L2_j_7_netPar1[19], dalpha_L2_j_7_netPar2[19] }), .SIGN({ SIGN_dalpha_L2_j_7_netPar0[19], SIGN_dalpha_L2_j_7_netPar1[19], SIGN_dalpha_L2_j_7_netPar2[19]}), .R_condition(rc[309]), .OUT(dalpha_L2_j_7[19]), .SIGN_out(SIGN_dalpha_L2_j_7[19]));
SS_ADDSUB ADDSUB_dalpha_L2_20_0(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_0_netPar0[20], dalpha_L2_j_0_netPar1[20], dalpha_L2_j_0_netPar2[20] }), .SIGN({ SIGN_dalpha_L2_j_0_netPar0[20], SIGN_dalpha_L2_j_0_netPar1[20], SIGN_dalpha_L2_j_0_netPar2[20]}), .R_condition(rc[310]), .OUT(dalpha_L2_j_0[20]), .SIGN_out(SIGN_dalpha_L2_j_0[20]));
SS_ADDSUB ADDSUB_dalpha_L2_20_1(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_1_netPar0[20], dalpha_L2_j_1_netPar1[20], dalpha_L2_j_1_netPar2[20] }), .SIGN({ SIGN_dalpha_L2_j_1_netPar0[20], SIGN_dalpha_L2_j_1_netPar1[20], SIGN_dalpha_L2_j_1_netPar2[20]}), .R_condition(rc[311]), .OUT(dalpha_L2_j_1[20]), .SIGN_out(SIGN_dalpha_L2_j_1[20]));
SS_ADDSUB ADDSUB_dalpha_L2_20_2(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_2_netPar0[20], dalpha_L2_j_2_netPar1[20], dalpha_L2_j_2_netPar2[20] }), .SIGN({ SIGN_dalpha_L2_j_2_netPar0[20], SIGN_dalpha_L2_j_2_netPar1[20], SIGN_dalpha_L2_j_2_netPar2[20]}), .R_condition(rc[312]), .OUT(dalpha_L2_j_2[20]), .SIGN_out(SIGN_dalpha_L2_j_2[20]));
SS_ADDSUB ADDSUB_dalpha_L2_20_3(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_3_netPar0[20], dalpha_L2_j_3_netPar1[20], dalpha_L2_j_3_netPar2[20] }), .SIGN({ SIGN_dalpha_L2_j_3_netPar0[20], SIGN_dalpha_L2_j_3_netPar1[20], SIGN_dalpha_L2_j_3_netPar2[20]}), .R_condition(rc[313]), .OUT(dalpha_L2_j_3[20]), .SIGN_out(SIGN_dalpha_L2_j_3[20]));
SS_ADDSUB ADDSUB_dalpha_L2_20_4(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_4_netPar0[20], dalpha_L2_j_4_netPar1[20], dalpha_L2_j_4_netPar2[20] }), .SIGN({ SIGN_dalpha_L2_j_4_netPar0[20], SIGN_dalpha_L2_j_4_netPar1[20], SIGN_dalpha_L2_j_4_netPar2[20]}), .R_condition(rc[314]), .OUT(dalpha_L2_j_4[20]), .SIGN_out(SIGN_dalpha_L2_j_4[20]));
SS_ADDSUB ADDSUB_dalpha_L2_20_5(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_5_netPar0[20], dalpha_L2_j_5_netPar1[20], dalpha_L2_j_5_netPar2[20] }), .SIGN({ SIGN_dalpha_L2_j_5_netPar0[20], SIGN_dalpha_L2_j_5_netPar1[20], SIGN_dalpha_L2_j_5_netPar2[20]}), .R_condition(rc[315]), .OUT(dalpha_L2_j_5[20]), .SIGN_out(SIGN_dalpha_L2_j_5[20]));
SS_ADDSUB ADDSUB_dalpha_L2_20_6(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_6_netPar0[20], dalpha_L2_j_6_netPar1[20], dalpha_L2_j_6_netPar2[20] }), .SIGN({ SIGN_dalpha_L2_j_6_netPar0[20], SIGN_dalpha_L2_j_6_netPar1[20], SIGN_dalpha_L2_j_6_netPar2[20]}), .R_condition(rc[316]), .OUT(dalpha_L2_j_6[20]), .SIGN_out(SIGN_dalpha_L2_j_6[20]));
SS_ADDSUB ADDSUB_dalpha_L2_20_7(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_7_netPar0[20], dalpha_L2_j_7_netPar1[20], dalpha_L2_j_7_netPar2[20] }), .SIGN({ SIGN_dalpha_L2_j_7_netPar0[20], SIGN_dalpha_L2_j_7_netPar1[20], SIGN_dalpha_L2_j_7_netPar2[20]}), .R_condition(rc[317]), .OUT(dalpha_L2_j_7[20]), .SIGN_out(SIGN_dalpha_L2_j_7[20]));
SS_ADDSUB ADDSUB_dalpha_L2_21_0(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_0_netPar0[21], dalpha_L2_j_0_netPar1[21], dalpha_L2_j_0_netPar2[21] }), .SIGN({ SIGN_dalpha_L2_j_0_netPar0[21], SIGN_dalpha_L2_j_0_netPar1[21], SIGN_dalpha_L2_j_0_netPar2[21]}), .R_condition(rc[318]), .OUT(dalpha_L2_j_0[21]), .SIGN_out(SIGN_dalpha_L2_j_0[21]));
SS_ADDSUB ADDSUB_dalpha_L2_21_1(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_1_netPar0[21], dalpha_L2_j_1_netPar1[21], dalpha_L2_j_1_netPar2[21] }), .SIGN({ SIGN_dalpha_L2_j_1_netPar0[21], SIGN_dalpha_L2_j_1_netPar1[21], SIGN_dalpha_L2_j_1_netPar2[21]}), .R_condition(rc[319]), .OUT(dalpha_L2_j_1[21]), .SIGN_out(SIGN_dalpha_L2_j_1[21]));
SS_ADDSUB ADDSUB_dalpha_L2_21_2(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_2_netPar0[21], dalpha_L2_j_2_netPar1[21], dalpha_L2_j_2_netPar2[21] }), .SIGN({ SIGN_dalpha_L2_j_2_netPar0[21], SIGN_dalpha_L2_j_2_netPar1[21], SIGN_dalpha_L2_j_2_netPar2[21]}), .R_condition(rc[320]), .OUT(dalpha_L2_j_2[21]), .SIGN_out(SIGN_dalpha_L2_j_2[21]));
SS_ADDSUB ADDSUB_dalpha_L2_21_3(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_3_netPar0[21], dalpha_L2_j_3_netPar1[21], dalpha_L2_j_3_netPar2[21] }), .SIGN({ SIGN_dalpha_L2_j_3_netPar0[21], SIGN_dalpha_L2_j_3_netPar1[21], SIGN_dalpha_L2_j_3_netPar2[21]}), .R_condition(rc[321]), .OUT(dalpha_L2_j_3[21]), .SIGN_out(SIGN_dalpha_L2_j_3[21]));
SS_ADDSUB ADDSUB_dalpha_L2_21_4(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_4_netPar0[21], dalpha_L2_j_4_netPar1[21], dalpha_L2_j_4_netPar2[21] }), .SIGN({ SIGN_dalpha_L2_j_4_netPar0[21], SIGN_dalpha_L2_j_4_netPar1[21], SIGN_dalpha_L2_j_4_netPar2[21]}), .R_condition(rc[322]), .OUT(dalpha_L2_j_4[21]), .SIGN_out(SIGN_dalpha_L2_j_4[21]));
SS_ADDSUB ADDSUB_dalpha_L2_21_5(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_5_netPar0[21], dalpha_L2_j_5_netPar1[21], dalpha_L2_j_5_netPar2[21] }), .SIGN({ SIGN_dalpha_L2_j_5_netPar0[21], SIGN_dalpha_L2_j_5_netPar1[21], SIGN_dalpha_L2_j_5_netPar2[21]}), .R_condition(rc[323]), .OUT(dalpha_L2_j_5[21]), .SIGN_out(SIGN_dalpha_L2_j_5[21]));
SS_ADDSUB ADDSUB_dalpha_L2_21_6(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_6_netPar0[21], dalpha_L2_j_6_netPar1[21], dalpha_L2_j_6_netPar2[21] }), .SIGN({ SIGN_dalpha_L2_j_6_netPar0[21], SIGN_dalpha_L2_j_6_netPar1[21], SIGN_dalpha_L2_j_6_netPar2[21]}), .R_condition(rc[324]), .OUT(dalpha_L2_j_6[21]), .SIGN_out(SIGN_dalpha_L2_j_6[21]));
SS_ADDSUB ADDSUB_dalpha_L2_21_7(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_7_netPar0[21], dalpha_L2_j_7_netPar1[21], dalpha_L2_j_7_netPar2[21] }), .SIGN({ SIGN_dalpha_L2_j_7_netPar0[21], SIGN_dalpha_L2_j_7_netPar1[21], SIGN_dalpha_L2_j_7_netPar2[21]}), .R_condition(rc[325]), .OUT(dalpha_L2_j_7[21]), .SIGN_out(SIGN_dalpha_L2_j_7[21]));
SS_ADDSUB ADDSUB_dalpha_L2_22_0(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_0_netPar0[22], dalpha_L2_j_0_netPar1[22], dalpha_L2_j_0_netPar2[22] }), .SIGN({ SIGN_dalpha_L2_j_0_netPar0[22], SIGN_dalpha_L2_j_0_netPar1[22], SIGN_dalpha_L2_j_0_netPar2[22]}), .R_condition(rc[326]), .OUT(dalpha_L2_j_0[22]), .SIGN_out(SIGN_dalpha_L2_j_0[22]));
SS_ADDSUB ADDSUB_dalpha_L2_22_1(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_1_netPar0[22], dalpha_L2_j_1_netPar1[22], dalpha_L2_j_1_netPar2[22] }), .SIGN({ SIGN_dalpha_L2_j_1_netPar0[22], SIGN_dalpha_L2_j_1_netPar1[22], SIGN_dalpha_L2_j_1_netPar2[22]}), .R_condition(rc[327]), .OUT(dalpha_L2_j_1[22]), .SIGN_out(SIGN_dalpha_L2_j_1[22]));
SS_ADDSUB ADDSUB_dalpha_L2_22_2(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_2_netPar0[22], dalpha_L2_j_2_netPar1[22], dalpha_L2_j_2_netPar2[22] }), .SIGN({ SIGN_dalpha_L2_j_2_netPar0[22], SIGN_dalpha_L2_j_2_netPar1[22], SIGN_dalpha_L2_j_2_netPar2[22]}), .R_condition(rc[328]), .OUT(dalpha_L2_j_2[22]), .SIGN_out(SIGN_dalpha_L2_j_2[22]));
SS_ADDSUB ADDSUB_dalpha_L2_22_3(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_3_netPar0[22], dalpha_L2_j_3_netPar1[22], dalpha_L2_j_3_netPar2[22] }), .SIGN({ SIGN_dalpha_L2_j_3_netPar0[22], SIGN_dalpha_L2_j_3_netPar1[22], SIGN_dalpha_L2_j_3_netPar2[22]}), .R_condition(rc[329]), .OUT(dalpha_L2_j_3[22]), .SIGN_out(SIGN_dalpha_L2_j_3[22]));
SS_ADDSUB ADDSUB_dalpha_L2_22_4(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_4_netPar0[22], dalpha_L2_j_4_netPar1[22], dalpha_L2_j_4_netPar2[22] }), .SIGN({ SIGN_dalpha_L2_j_4_netPar0[22], SIGN_dalpha_L2_j_4_netPar1[22], SIGN_dalpha_L2_j_4_netPar2[22]}), .R_condition(rc[330]), .OUT(dalpha_L2_j_4[22]), .SIGN_out(SIGN_dalpha_L2_j_4[22]));
SS_ADDSUB ADDSUB_dalpha_L2_22_5(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_5_netPar0[22], dalpha_L2_j_5_netPar1[22], dalpha_L2_j_5_netPar2[22] }), .SIGN({ SIGN_dalpha_L2_j_5_netPar0[22], SIGN_dalpha_L2_j_5_netPar1[22], SIGN_dalpha_L2_j_5_netPar2[22]}), .R_condition(rc[331]), .OUT(dalpha_L2_j_5[22]), .SIGN_out(SIGN_dalpha_L2_j_5[22]));
SS_ADDSUB ADDSUB_dalpha_L2_22_6(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_6_netPar0[22], dalpha_L2_j_6_netPar1[22], dalpha_L2_j_6_netPar2[22] }), .SIGN({ SIGN_dalpha_L2_j_6_netPar0[22], SIGN_dalpha_L2_j_6_netPar1[22], SIGN_dalpha_L2_j_6_netPar2[22]}), .R_condition(rc[332]), .OUT(dalpha_L2_j_6[22]), .SIGN_out(SIGN_dalpha_L2_j_6[22]));
SS_ADDSUB ADDSUB_dalpha_L2_22_7(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_7_netPar0[22], dalpha_L2_j_7_netPar1[22], dalpha_L2_j_7_netPar2[22] }), .SIGN({ SIGN_dalpha_L2_j_7_netPar0[22], SIGN_dalpha_L2_j_7_netPar1[22], SIGN_dalpha_L2_j_7_netPar2[22]}), .R_condition(rc[333]), .OUT(dalpha_L2_j_7[22]), .SIGN_out(SIGN_dalpha_L2_j_7[22]));
SS_ADDSUB ADDSUB_dalpha_L2_23_0(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_0_netPar0[23], dalpha_L2_j_0_netPar1[23], dalpha_L2_j_0_netPar2[23] }), .SIGN({ SIGN_dalpha_L2_j_0_netPar0[23], SIGN_dalpha_L2_j_0_netPar1[23], SIGN_dalpha_L2_j_0_netPar2[23]}), .R_condition(rc[334]), .OUT(dalpha_L2_j_0[23]), .SIGN_out(SIGN_dalpha_L2_j_0[23]));
SS_ADDSUB ADDSUB_dalpha_L2_23_1(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_1_netPar0[23], dalpha_L2_j_1_netPar1[23], dalpha_L2_j_1_netPar2[23] }), .SIGN({ SIGN_dalpha_L2_j_1_netPar0[23], SIGN_dalpha_L2_j_1_netPar1[23], SIGN_dalpha_L2_j_1_netPar2[23]}), .R_condition(rc[335]), .OUT(dalpha_L2_j_1[23]), .SIGN_out(SIGN_dalpha_L2_j_1[23]));
SS_ADDSUB ADDSUB_dalpha_L2_23_2(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_2_netPar0[23], dalpha_L2_j_2_netPar1[23], dalpha_L2_j_2_netPar2[23] }), .SIGN({ SIGN_dalpha_L2_j_2_netPar0[23], SIGN_dalpha_L2_j_2_netPar1[23], SIGN_dalpha_L2_j_2_netPar2[23]}), .R_condition(rc[336]), .OUT(dalpha_L2_j_2[23]), .SIGN_out(SIGN_dalpha_L2_j_2[23]));
SS_ADDSUB ADDSUB_dalpha_L2_23_3(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_3_netPar0[23], dalpha_L2_j_3_netPar1[23], dalpha_L2_j_3_netPar2[23] }), .SIGN({ SIGN_dalpha_L2_j_3_netPar0[23], SIGN_dalpha_L2_j_3_netPar1[23], SIGN_dalpha_L2_j_3_netPar2[23]}), .R_condition(rc[337]), .OUT(dalpha_L2_j_3[23]), .SIGN_out(SIGN_dalpha_L2_j_3[23]));
SS_ADDSUB ADDSUB_dalpha_L2_23_4(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_4_netPar0[23], dalpha_L2_j_4_netPar1[23], dalpha_L2_j_4_netPar2[23] }), .SIGN({ SIGN_dalpha_L2_j_4_netPar0[23], SIGN_dalpha_L2_j_4_netPar1[23], SIGN_dalpha_L2_j_4_netPar2[23]}), .R_condition(rc[338]), .OUT(dalpha_L2_j_4[23]), .SIGN_out(SIGN_dalpha_L2_j_4[23]));
SS_ADDSUB ADDSUB_dalpha_L2_23_5(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_5_netPar0[23], dalpha_L2_j_5_netPar1[23], dalpha_L2_j_5_netPar2[23] }), .SIGN({ SIGN_dalpha_L2_j_5_netPar0[23], SIGN_dalpha_L2_j_5_netPar1[23], SIGN_dalpha_L2_j_5_netPar2[23]}), .R_condition(rc[339]), .OUT(dalpha_L2_j_5[23]), .SIGN_out(SIGN_dalpha_L2_j_5[23]));
SS_ADDSUB ADDSUB_dalpha_L2_23_6(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_6_netPar0[23], dalpha_L2_j_6_netPar1[23], dalpha_L2_j_6_netPar2[23] }), .SIGN({ SIGN_dalpha_L2_j_6_netPar0[23], SIGN_dalpha_L2_j_6_netPar1[23], SIGN_dalpha_L2_j_6_netPar2[23]}), .R_condition(rc[340]), .OUT(dalpha_L2_j_6[23]), .SIGN_out(SIGN_dalpha_L2_j_6[23]));
SS_ADDSUB ADDSUB_dalpha_L2_23_7(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_7_netPar0[23], dalpha_L2_j_7_netPar1[23], dalpha_L2_j_7_netPar2[23] }), .SIGN({ SIGN_dalpha_L2_j_7_netPar0[23], SIGN_dalpha_L2_j_7_netPar1[23], SIGN_dalpha_L2_j_7_netPar2[23]}), .R_condition(rc[341]), .OUT(dalpha_L2_j_7[23]), .SIGN_out(SIGN_dalpha_L2_j_7[23]));
SS_ADDSUB ADDSUB_dalpha_L2_24_0(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_0_netPar0[24], dalpha_L2_j_0_netPar1[24], dalpha_L2_j_0_netPar2[24] }), .SIGN({ SIGN_dalpha_L2_j_0_netPar0[24], SIGN_dalpha_L2_j_0_netPar1[24], SIGN_dalpha_L2_j_0_netPar2[24]}), .R_condition(rc[342]), .OUT(dalpha_L2_j_0[24]), .SIGN_out(SIGN_dalpha_L2_j_0[24]));
SS_ADDSUB ADDSUB_dalpha_L2_24_1(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_1_netPar0[24], dalpha_L2_j_1_netPar1[24], dalpha_L2_j_1_netPar2[24] }), .SIGN({ SIGN_dalpha_L2_j_1_netPar0[24], SIGN_dalpha_L2_j_1_netPar1[24], SIGN_dalpha_L2_j_1_netPar2[24]}), .R_condition(rc[343]), .OUT(dalpha_L2_j_1[24]), .SIGN_out(SIGN_dalpha_L2_j_1[24]));
SS_ADDSUB ADDSUB_dalpha_L2_24_2(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_2_netPar0[24], dalpha_L2_j_2_netPar1[24], dalpha_L2_j_2_netPar2[24] }), .SIGN({ SIGN_dalpha_L2_j_2_netPar0[24], SIGN_dalpha_L2_j_2_netPar1[24], SIGN_dalpha_L2_j_2_netPar2[24]}), .R_condition(rc[344]), .OUT(dalpha_L2_j_2[24]), .SIGN_out(SIGN_dalpha_L2_j_2[24]));
SS_ADDSUB ADDSUB_dalpha_L2_24_3(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_3_netPar0[24], dalpha_L2_j_3_netPar1[24], dalpha_L2_j_3_netPar2[24] }), .SIGN({ SIGN_dalpha_L2_j_3_netPar0[24], SIGN_dalpha_L2_j_3_netPar1[24], SIGN_dalpha_L2_j_3_netPar2[24]}), .R_condition(rc[345]), .OUT(dalpha_L2_j_3[24]), .SIGN_out(SIGN_dalpha_L2_j_3[24]));
SS_ADDSUB ADDSUB_dalpha_L2_24_4(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_4_netPar0[24], dalpha_L2_j_4_netPar1[24], dalpha_L2_j_4_netPar2[24] }), .SIGN({ SIGN_dalpha_L2_j_4_netPar0[24], SIGN_dalpha_L2_j_4_netPar1[24], SIGN_dalpha_L2_j_4_netPar2[24]}), .R_condition(rc[346]), .OUT(dalpha_L2_j_4[24]), .SIGN_out(SIGN_dalpha_L2_j_4[24]));
SS_ADDSUB ADDSUB_dalpha_L2_24_5(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_5_netPar0[24], dalpha_L2_j_5_netPar1[24], dalpha_L2_j_5_netPar2[24] }), .SIGN({ SIGN_dalpha_L2_j_5_netPar0[24], SIGN_dalpha_L2_j_5_netPar1[24], SIGN_dalpha_L2_j_5_netPar2[24]}), .R_condition(rc[347]), .OUT(dalpha_L2_j_5[24]), .SIGN_out(SIGN_dalpha_L2_j_5[24]));
SS_ADDSUB ADDSUB_dalpha_L2_24_6(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_6_netPar0[24], dalpha_L2_j_6_netPar1[24], dalpha_L2_j_6_netPar2[24] }), .SIGN({ SIGN_dalpha_L2_j_6_netPar0[24], SIGN_dalpha_L2_j_6_netPar1[24], SIGN_dalpha_L2_j_6_netPar2[24]}), .R_condition(rc[348]), .OUT(dalpha_L2_j_6[24]), .SIGN_out(SIGN_dalpha_L2_j_6[24]));
SS_ADDSUB ADDSUB_dalpha_L2_24_7(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L2_j_7_netPar0[24], dalpha_L2_j_7_netPar1[24], dalpha_L2_j_7_netPar2[24] }), .SIGN({ SIGN_dalpha_L2_j_7_netPar0[24], SIGN_dalpha_L2_j_7_netPar1[24], SIGN_dalpha_L2_j_7_netPar2[24]}), .R_condition(rc[349]), .OUT(dalpha_L2_j_7[24]), .SIGN_out(SIGN_dalpha_L2_j_7[24]));
defparam ADDSUB_dalpha_L2_0_0.N = 3;
defparam ADDSUB_dalpha_L2_0_1.N = 3;
defparam ADDSUB_dalpha_L2_0_2.N = 3;
defparam ADDSUB_dalpha_L2_0_3.N = 3;
defparam ADDSUB_dalpha_L2_0_4.N = 3;
defparam ADDSUB_dalpha_L2_0_5.N = 3;
defparam ADDSUB_dalpha_L2_0_6.N = 3;
defparam ADDSUB_dalpha_L2_0_7.N = 3;
defparam ADDSUB_dalpha_L2_1_0.N = 3;
defparam ADDSUB_dalpha_L2_1_1.N = 3;
defparam ADDSUB_dalpha_L2_1_2.N = 3;
defparam ADDSUB_dalpha_L2_1_3.N = 3;
defparam ADDSUB_dalpha_L2_1_4.N = 3;
defparam ADDSUB_dalpha_L2_1_5.N = 3;
defparam ADDSUB_dalpha_L2_1_6.N = 3;
defparam ADDSUB_dalpha_L2_1_7.N = 3;
defparam ADDSUB_dalpha_L2_2_0.N = 3;
defparam ADDSUB_dalpha_L2_2_1.N = 3;
defparam ADDSUB_dalpha_L2_2_2.N = 3;
defparam ADDSUB_dalpha_L2_2_3.N = 3;
defparam ADDSUB_dalpha_L2_2_4.N = 3;
defparam ADDSUB_dalpha_L2_2_5.N = 3;
defparam ADDSUB_dalpha_L2_2_6.N = 3;
defparam ADDSUB_dalpha_L2_2_7.N = 3;
defparam ADDSUB_dalpha_L2_3_0.N = 3;
defparam ADDSUB_dalpha_L2_3_1.N = 3;
defparam ADDSUB_dalpha_L2_3_2.N = 3;
defparam ADDSUB_dalpha_L2_3_3.N = 3;
defparam ADDSUB_dalpha_L2_3_4.N = 3;
defparam ADDSUB_dalpha_L2_3_5.N = 3;
defparam ADDSUB_dalpha_L2_3_6.N = 3;
defparam ADDSUB_dalpha_L2_3_7.N = 3;
defparam ADDSUB_dalpha_L2_4_0.N = 3;
defparam ADDSUB_dalpha_L2_4_1.N = 3;
defparam ADDSUB_dalpha_L2_4_2.N = 3;
defparam ADDSUB_dalpha_L2_4_3.N = 3;
defparam ADDSUB_dalpha_L2_4_4.N = 3;
defparam ADDSUB_dalpha_L2_4_5.N = 3;
defparam ADDSUB_dalpha_L2_4_6.N = 3;
defparam ADDSUB_dalpha_L2_4_7.N = 3;
defparam ADDSUB_dalpha_L2_5_0.N = 3;
defparam ADDSUB_dalpha_L2_5_1.N = 3;
defparam ADDSUB_dalpha_L2_5_2.N = 3;
defparam ADDSUB_dalpha_L2_5_3.N = 3;
defparam ADDSUB_dalpha_L2_5_4.N = 3;
defparam ADDSUB_dalpha_L2_5_5.N = 3;
defparam ADDSUB_dalpha_L2_5_6.N = 3;
defparam ADDSUB_dalpha_L2_5_7.N = 3;
defparam ADDSUB_dalpha_L2_6_0.N = 3;
defparam ADDSUB_dalpha_L2_6_1.N = 3;
defparam ADDSUB_dalpha_L2_6_2.N = 3;
defparam ADDSUB_dalpha_L2_6_3.N = 3;
defparam ADDSUB_dalpha_L2_6_4.N = 3;
defparam ADDSUB_dalpha_L2_6_5.N = 3;
defparam ADDSUB_dalpha_L2_6_6.N = 3;
defparam ADDSUB_dalpha_L2_6_7.N = 3;
defparam ADDSUB_dalpha_L2_7_0.N = 3;
defparam ADDSUB_dalpha_L2_7_1.N = 3;
defparam ADDSUB_dalpha_L2_7_2.N = 3;
defparam ADDSUB_dalpha_L2_7_3.N = 3;
defparam ADDSUB_dalpha_L2_7_4.N = 3;
defparam ADDSUB_dalpha_L2_7_5.N = 3;
defparam ADDSUB_dalpha_L2_7_6.N = 3;
defparam ADDSUB_dalpha_L2_7_7.N = 3;
defparam ADDSUB_dalpha_L2_8_0.N = 3;
defparam ADDSUB_dalpha_L2_8_1.N = 3;
defparam ADDSUB_dalpha_L2_8_2.N = 3;
defparam ADDSUB_dalpha_L2_8_3.N = 3;
defparam ADDSUB_dalpha_L2_8_4.N = 3;
defparam ADDSUB_dalpha_L2_8_5.N = 3;
defparam ADDSUB_dalpha_L2_8_6.N = 3;
defparam ADDSUB_dalpha_L2_8_7.N = 3;
defparam ADDSUB_dalpha_L2_9_0.N = 3;
defparam ADDSUB_dalpha_L2_9_1.N = 3;
defparam ADDSUB_dalpha_L2_9_2.N = 3;
defparam ADDSUB_dalpha_L2_9_3.N = 3;
defparam ADDSUB_dalpha_L2_9_4.N = 3;
defparam ADDSUB_dalpha_L2_9_5.N = 3;
defparam ADDSUB_dalpha_L2_9_6.N = 3;
defparam ADDSUB_dalpha_L2_9_7.N = 3;
defparam ADDSUB_dalpha_L2_10_0.N = 3;
defparam ADDSUB_dalpha_L2_10_1.N = 3;
defparam ADDSUB_dalpha_L2_10_2.N = 3;
defparam ADDSUB_dalpha_L2_10_3.N = 3;
defparam ADDSUB_dalpha_L2_10_4.N = 3;
defparam ADDSUB_dalpha_L2_10_5.N = 3;
defparam ADDSUB_dalpha_L2_10_6.N = 3;
defparam ADDSUB_dalpha_L2_10_7.N = 3;
defparam ADDSUB_dalpha_L2_11_0.N = 3;
defparam ADDSUB_dalpha_L2_11_1.N = 3;
defparam ADDSUB_dalpha_L2_11_2.N = 3;
defparam ADDSUB_dalpha_L2_11_3.N = 3;
defparam ADDSUB_dalpha_L2_11_4.N = 3;
defparam ADDSUB_dalpha_L2_11_5.N = 3;
defparam ADDSUB_dalpha_L2_11_6.N = 3;
defparam ADDSUB_dalpha_L2_11_7.N = 3;
defparam ADDSUB_dalpha_L2_12_0.N = 3;
defparam ADDSUB_dalpha_L2_12_1.N = 3;
defparam ADDSUB_dalpha_L2_12_2.N = 3;
defparam ADDSUB_dalpha_L2_12_3.N = 3;
defparam ADDSUB_dalpha_L2_12_4.N = 3;
defparam ADDSUB_dalpha_L2_12_5.N = 3;
defparam ADDSUB_dalpha_L2_12_6.N = 3;
defparam ADDSUB_dalpha_L2_12_7.N = 3;
defparam ADDSUB_dalpha_L2_13_0.N = 3;
defparam ADDSUB_dalpha_L2_13_1.N = 3;
defparam ADDSUB_dalpha_L2_13_2.N = 3;
defparam ADDSUB_dalpha_L2_13_3.N = 3;
defparam ADDSUB_dalpha_L2_13_4.N = 3;
defparam ADDSUB_dalpha_L2_13_5.N = 3;
defparam ADDSUB_dalpha_L2_13_6.N = 3;
defparam ADDSUB_dalpha_L2_13_7.N = 3;
defparam ADDSUB_dalpha_L2_14_0.N = 3;
defparam ADDSUB_dalpha_L2_14_1.N = 3;
defparam ADDSUB_dalpha_L2_14_2.N = 3;
defparam ADDSUB_dalpha_L2_14_3.N = 3;
defparam ADDSUB_dalpha_L2_14_4.N = 3;
defparam ADDSUB_dalpha_L2_14_5.N = 3;
defparam ADDSUB_dalpha_L2_14_6.N = 3;
defparam ADDSUB_dalpha_L2_14_7.N = 3;
defparam ADDSUB_dalpha_L2_15_0.N = 3;
defparam ADDSUB_dalpha_L2_15_1.N = 3;
defparam ADDSUB_dalpha_L2_15_2.N = 3;
defparam ADDSUB_dalpha_L2_15_3.N = 3;
defparam ADDSUB_dalpha_L2_15_4.N = 3;
defparam ADDSUB_dalpha_L2_15_5.N = 3;
defparam ADDSUB_dalpha_L2_15_6.N = 3;
defparam ADDSUB_dalpha_L2_15_7.N = 3;
defparam ADDSUB_dalpha_L2_16_0.N = 3;
defparam ADDSUB_dalpha_L2_16_1.N = 3;
defparam ADDSUB_dalpha_L2_16_2.N = 3;
defparam ADDSUB_dalpha_L2_16_3.N = 3;
defparam ADDSUB_dalpha_L2_16_4.N = 3;
defparam ADDSUB_dalpha_L2_16_5.N = 3;
defparam ADDSUB_dalpha_L2_16_6.N = 3;
defparam ADDSUB_dalpha_L2_16_7.N = 3;
defparam ADDSUB_dalpha_L2_17_0.N = 3;
defparam ADDSUB_dalpha_L2_17_1.N = 3;
defparam ADDSUB_dalpha_L2_17_2.N = 3;
defparam ADDSUB_dalpha_L2_17_3.N = 3;
defparam ADDSUB_dalpha_L2_17_4.N = 3;
defparam ADDSUB_dalpha_L2_17_5.N = 3;
defparam ADDSUB_dalpha_L2_17_6.N = 3;
defparam ADDSUB_dalpha_L2_17_7.N = 3;
defparam ADDSUB_dalpha_L2_18_0.N = 3;
defparam ADDSUB_dalpha_L2_18_1.N = 3;
defparam ADDSUB_dalpha_L2_18_2.N = 3;
defparam ADDSUB_dalpha_L2_18_3.N = 3;
defparam ADDSUB_dalpha_L2_18_4.N = 3;
defparam ADDSUB_dalpha_L2_18_5.N = 3;
defparam ADDSUB_dalpha_L2_18_6.N = 3;
defparam ADDSUB_dalpha_L2_18_7.N = 3;
defparam ADDSUB_dalpha_L2_19_0.N = 3;
defparam ADDSUB_dalpha_L2_19_1.N = 3;
defparam ADDSUB_dalpha_L2_19_2.N = 3;
defparam ADDSUB_dalpha_L2_19_3.N = 3;
defparam ADDSUB_dalpha_L2_19_4.N = 3;
defparam ADDSUB_dalpha_L2_19_5.N = 3;
defparam ADDSUB_dalpha_L2_19_6.N = 3;
defparam ADDSUB_dalpha_L2_19_7.N = 3;
defparam ADDSUB_dalpha_L2_20_0.N = 3;
defparam ADDSUB_dalpha_L2_20_1.N = 3;
defparam ADDSUB_dalpha_L2_20_2.N = 3;
defparam ADDSUB_dalpha_L2_20_3.N = 3;
defparam ADDSUB_dalpha_L2_20_4.N = 3;
defparam ADDSUB_dalpha_L2_20_5.N = 3;
defparam ADDSUB_dalpha_L2_20_6.N = 3;
defparam ADDSUB_dalpha_L2_20_7.N = 3;
defparam ADDSUB_dalpha_L2_21_0.N = 3;
defparam ADDSUB_dalpha_L2_21_1.N = 3;
defparam ADDSUB_dalpha_L2_21_2.N = 3;
defparam ADDSUB_dalpha_L2_21_3.N = 3;
defparam ADDSUB_dalpha_L2_21_4.N = 3;
defparam ADDSUB_dalpha_L2_21_5.N = 3;
defparam ADDSUB_dalpha_L2_21_6.N = 3;
defparam ADDSUB_dalpha_L2_21_7.N = 3;
defparam ADDSUB_dalpha_L2_22_0.N = 3;
defparam ADDSUB_dalpha_L2_22_1.N = 3;
defparam ADDSUB_dalpha_L2_22_2.N = 3;
defparam ADDSUB_dalpha_L2_22_3.N = 3;
defparam ADDSUB_dalpha_L2_22_4.N = 3;
defparam ADDSUB_dalpha_L2_22_5.N = 3;
defparam ADDSUB_dalpha_L2_22_6.N = 3;
defparam ADDSUB_dalpha_L2_22_7.N = 3;
defparam ADDSUB_dalpha_L2_23_0.N = 3;
defparam ADDSUB_dalpha_L2_23_1.N = 3;
defparam ADDSUB_dalpha_L2_23_2.N = 3;
defparam ADDSUB_dalpha_L2_23_3.N = 3;
defparam ADDSUB_dalpha_L2_23_4.N = 3;
defparam ADDSUB_dalpha_L2_23_5.N = 3;
defparam ADDSUB_dalpha_L2_23_6.N = 3;
defparam ADDSUB_dalpha_L2_23_7.N = 3;
defparam ADDSUB_dalpha_L2_24_0.N = 3;
defparam ADDSUB_dalpha_L2_24_1.N = 3;
defparam ADDSUB_dalpha_L2_24_2.N = 3;
defparam ADDSUB_dalpha_L2_24_3.N = 3;
defparam ADDSUB_dalpha_L2_24_4.N = 3;
defparam ADDSUB_dalpha_L2_24_5.N = 3;
defparam ADDSUB_dalpha_L2_24_6.N = 3;
defparam ADDSUB_dalpha_L2_24_7.N = 3;
defparam ADDSUB_dalpha_L2_0_0.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_0_1.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_0_2.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_0_3.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_0_4.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_0_5.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_0_6.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_0_7.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_1_0.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_1_1.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_1_2.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_1_3.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_1_4.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_1_5.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_1_6.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_1_7.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_2_0.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_2_1.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_2_2.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_2_3.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_2_4.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_2_5.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_2_6.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_2_7.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_3_0.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_3_1.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_3_2.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_3_3.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_3_4.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_3_5.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_3_6.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_3_7.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_4_0.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_4_1.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_4_2.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_4_3.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_4_4.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_4_5.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_4_6.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_4_7.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_5_0.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_5_1.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_5_2.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_5_3.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_5_4.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_5_5.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_5_6.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_5_7.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_6_0.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_6_1.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_6_2.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_6_3.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_6_4.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_6_5.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_6_6.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_6_7.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_7_0.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_7_1.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_7_2.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_7_3.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_7_4.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_7_5.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_7_6.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_7_7.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_8_0.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_8_1.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_8_2.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_8_3.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_8_4.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_8_5.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_8_6.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_8_7.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_9_0.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_9_1.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_9_2.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_9_3.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_9_4.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_9_5.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_9_6.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_9_7.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_10_0.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_10_1.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_10_2.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_10_3.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_10_4.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_10_5.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_10_6.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_10_7.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_11_0.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_11_1.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_11_2.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_11_3.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_11_4.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_11_5.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_11_6.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_11_7.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_12_0.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_12_1.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_12_2.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_12_3.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_12_4.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_12_5.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_12_6.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_12_7.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_13_0.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_13_1.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_13_2.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_13_3.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_13_4.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_13_5.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_13_6.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_13_7.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_14_0.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_14_1.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_14_2.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_14_3.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_14_4.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_14_5.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_14_6.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_14_7.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_15_0.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_15_1.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_15_2.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_15_3.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_15_4.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_15_5.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_15_6.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_15_7.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_16_0.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_16_1.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_16_2.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_16_3.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_16_4.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_16_5.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_16_6.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_16_7.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_17_0.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_17_1.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_17_2.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_17_3.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_17_4.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_17_5.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_17_6.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_17_7.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_18_0.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_18_1.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_18_2.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_18_3.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_18_4.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_18_5.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_18_6.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_18_7.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_19_0.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_19_1.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_19_2.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_19_3.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_19_4.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_19_5.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_19_6.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_19_7.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_20_0.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_20_1.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_20_2.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_20_3.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_20_4.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_20_5.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_20_6.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_20_7.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_21_0.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_21_1.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_21_2.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_21_3.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_21_4.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_21_5.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_21_6.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_21_7.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_22_0.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_22_1.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_22_2.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_22_3.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_22_4.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_22_5.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_22_6.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_22_7.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_23_0.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_23_1.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_23_2.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_23_3.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_23_4.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_23_5.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_23_6.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_23_7.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_24_0.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_24_1.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_24_2.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_24_3.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_24_4.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_24_5.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_24_6.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L2_24_7.DIFFCOUNTER_SIZE = 3;

SS_ADDSUB ADDSUB_dbeta_L2_0(.CLK(CLK), .INIT(INIT), .IN({ dbeta_L2_netPar0[0], dbeta_L2_netPar1[0], dbeta_L2_netPar2[0] }), .SIGN({ SIGN_dbeta_L2_netPar0[0], SIGN_dbeta_L2_netPar1[0], SIGN_dbeta_L2_netPar2[0]}), .R_condition(rc[350]), .OUT(dbeta_L2[0]), .SIGN_out(SIGN_dbeta_L2[0]));
SS_ADDSUB ADDSUB_dbeta_L2_1(.CLK(CLK), .INIT(INIT), .IN({ dbeta_L2_netPar0[1], dbeta_L2_netPar1[1], dbeta_L2_netPar2[1] }), .SIGN({ SIGN_dbeta_L2_netPar0[1], SIGN_dbeta_L2_netPar1[1], SIGN_dbeta_L2_netPar2[1]}), .R_condition(rc[351]), .OUT(dbeta_L2[1]), .SIGN_out(SIGN_dbeta_L2[1]));
SS_ADDSUB ADDSUB_dbeta_L2_2(.CLK(CLK), .INIT(INIT), .IN({ dbeta_L2_netPar0[2], dbeta_L2_netPar1[2], dbeta_L2_netPar2[2] }), .SIGN({ SIGN_dbeta_L2_netPar0[2], SIGN_dbeta_L2_netPar1[2], SIGN_dbeta_L2_netPar2[2]}), .R_condition(rc[352]), .OUT(dbeta_L2[2]), .SIGN_out(SIGN_dbeta_L2[2]));
SS_ADDSUB ADDSUB_dbeta_L2_3(.CLK(CLK), .INIT(INIT), .IN({ dbeta_L2_netPar0[3], dbeta_L2_netPar1[3], dbeta_L2_netPar2[3] }), .SIGN({ SIGN_dbeta_L2_netPar0[3], SIGN_dbeta_L2_netPar1[3], SIGN_dbeta_L2_netPar2[3]}), .R_condition(rc[353]), .OUT(dbeta_L2[3]), .SIGN_out(SIGN_dbeta_L2[3]));
SS_ADDSUB ADDSUB_dbeta_L2_4(.CLK(CLK), .INIT(INIT), .IN({ dbeta_L2_netPar0[4], dbeta_L2_netPar1[4], dbeta_L2_netPar2[4] }), .SIGN({ SIGN_dbeta_L2_netPar0[4], SIGN_dbeta_L2_netPar1[4], SIGN_dbeta_L2_netPar2[4]}), .R_condition(rc[354]), .OUT(dbeta_L2[4]), .SIGN_out(SIGN_dbeta_L2[4]));
SS_ADDSUB ADDSUB_dbeta_L2_5(.CLK(CLK), .INIT(INIT), .IN({ dbeta_L2_netPar0[5], dbeta_L2_netPar1[5], dbeta_L2_netPar2[5] }), .SIGN({ SIGN_dbeta_L2_netPar0[5], SIGN_dbeta_L2_netPar1[5], SIGN_dbeta_L2_netPar2[5]}), .R_condition(rc[355]), .OUT(dbeta_L2[5]), .SIGN_out(SIGN_dbeta_L2[5]));
SS_ADDSUB ADDSUB_dbeta_L2_6(.CLK(CLK), .INIT(INIT), .IN({ dbeta_L2_netPar0[6], dbeta_L2_netPar1[6], dbeta_L2_netPar2[6] }), .SIGN({ SIGN_dbeta_L2_netPar0[6], SIGN_dbeta_L2_netPar1[6], SIGN_dbeta_L2_netPar2[6]}), .R_condition(rc[356]), .OUT(dbeta_L2[6]), .SIGN_out(SIGN_dbeta_L2[6]));
SS_ADDSUB ADDSUB_dbeta_L2_7(.CLK(CLK), .INIT(INIT), .IN({ dbeta_L2_netPar0[7], dbeta_L2_netPar1[7], dbeta_L2_netPar2[7] }), .SIGN({ SIGN_dbeta_L2_netPar0[7], SIGN_dbeta_L2_netPar1[7], SIGN_dbeta_L2_netPar2[7]}), .R_condition(rc[357]), .OUT(dbeta_L2[7]), .SIGN_out(SIGN_dbeta_L2[7]));
defparam ADDSUB_dbeta_L2_0.N = 3;
defparam ADDSUB_dbeta_L2_1.N = 3;
defparam ADDSUB_dbeta_L2_2.N = 3;
defparam ADDSUB_dbeta_L2_3.N = 3;
defparam ADDSUB_dbeta_L2_4.N = 3;
defparam ADDSUB_dbeta_L2_5.N = 3;
defparam ADDSUB_dbeta_L2_6.N = 3;
defparam ADDSUB_dbeta_L2_7.N = 3;
defparam ADDSUB_dbeta_L2_0.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dbeta_L2_1.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dbeta_L2_2.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dbeta_L2_3.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dbeta_L2_4.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dbeta_L2_5.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dbeta_L2_6.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dbeta_L2_7.DIFFCOUNTER_SIZE = 3;


SS_ADDSUB ADDSUB_dalpha_L3_0_0(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L3_j_0_netPar0[0], dalpha_L3_j_0_netPar1[0], dalpha_L3_j_0_netPar2[0] }), .SIGN({ SIGN_dalpha_L3_j_0_netPar0[0], SIGN_dalpha_L3_j_0_netPar1[0], SIGN_dalpha_L3_j_0_netPar2[0]}), .R_condition(rc[358]), .OUT(dalpha_L3_j_0[0]), .SIGN_out(SIGN_dalpha_L3_j_0[0]));
SS_ADDSUB ADDSUB_dalpha_L3_0_1(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L3_j_1_netPar0[0], dalpha_L3_j_1_netPar1[0], dalpha_L3_j_1_netPar2[0] }), .SIGN({ SIGN_dalpha_L3_j_1_netPar0[0], SIGN_dalpha_L3_j_1_netPar1[0], SIGN_dalpha_L3_j_1_netPar2[0]}), .R_condition(rc[359]), .OUT(dalpha_L3_j_1[0]), .SIGN_out(SIGN_dalpha_L3_j_1[0]));
SS_ADDSUB ADDSUB_dalpha_L3_0_2(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L3_j_2_netPar0[0], dalpha_L3_j_2_netPar1[0], dalpha_L3_j_2_netPar2[0] }), .SIGN({ SIGN_dalpha_L3_j_2_netPar0[0], SIGN_dalpha_L3_j_2_netPar1[0], SIGN_dalpha_L3_j_2_netPar2[0]}), .R_condition(rc[360]), .OUT(dalpha_L3_j_2[0]), .SIGN_out(SIGN_dalpha_L3_j_2[0]));
SS_ADDSUB ADDSUB_dalpha_L3_0_3(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L3_j_3_netPar0[0], dalpha_L3_j_3_netPar1[0], dalpha_L3_j_3_netPar2[0] }), .SIGN({ SIGN_dalpha_L3_j_3_netPar0[0], SIGN_dalpha_L3_j_3_netPar1[0], SIGN_dalpha_L3_j_3_netPar2[0]}), .R_condition(rc[361]), .OUT(dalpha_L3_j_3[0]), .SIGN_out(SIGN_dalpha_L3_j_3[0]));
SS_ADDSUB ADDSUB_dalpha_L3_0_4(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L3_j_4_netPar0[0], dalpha_L3_j_4_netPar1[0], dalpha_L3_j_4_netPar2[0] }), .SIGN({ SIGN_dalpha_L3_j_4_netPar0[0], SIGN_dalpha_L3_j_4_netPar1[0], SIGN_dalpha_L3_j_4_netPar2[0]}), .R_condition(rc[362]), .OUT(dalpha_L3_j_4[0]), .SIGN_out(SIGN_dalpha_L3_j_4[0]));
SS_ADDSUB ADDSUB_dalpha_L3_1_0(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L3_j_0_netPar0[1], dalpha_L3_j_0_netPar1[1], dalpha_L3_j_0_netPar2[1] }), .SIGN({ SIGN_dalpha_L3_j_0_netPar0[1], SIGN_dalpha_L3_j_0_netPar1[1], SIGN_dalpha_L3_j_0_netPar2[1]}), .R_condition(rc[363]), .OUT(dalpha_L3_j_0[1]), .SIGN_out(SIGN_dalpha_L3_j_0[1]));
SS_ADDSUB ADDSUB_dalpha_L3_1_1(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L3_j_1_netPar0[1], dalpha_L3_j_1_netPar1[1], dalpha_L3_j_1_netPar2[1] }), .SIGN({ SIGN_dalpha_L3_j_1_netPar0[1], SIGN_dalpha_L3_j_1_netPar1[1], SIGN_dalpha_L3_j_1_netPar2[1]}), .R_condition(rc[364]), .OUT(dalpha_L3_j_1[1]), .SIGN_out(SIGN_dalpha_L3_j_1[1]));
SS_ADDSUB ADDSUB_dalpha_L3_1_2(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L3_j_2_netPar0[1], dalpha_L3_j_2_netPar1[1], dalpha_L3_j_2_netPar2[1] }), .SIGN({ SIGN_dalpha_L3_j_2_netPar0[1], SIGN_dalpha_L3_j_2_netPar1[1], SIGN_dalpha_L3_j_2_netPar2[1]}), .R_condition(rc[365]), .OUT(dalpha_L3_j_2[1]), .SIGN_out(SIGN_dalpha_L3_j_2[1]));
SS_ADDSUB ADDSUB_dalpha_L3_1_3(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L3_j_3_netPar0[1], dalpha_L3_j_3_netPar1[1], dalpha_L3_j_3_netPar2[1] }), .SIGN({ SIGN_dalpha_L3_j_3_netPar0[1], SIGN_dalpha_L3_j_3_netPar1[1], SIGN_dalpha_L3_j_3_netPar2[1]}), .R_condition(rc[366]), .OUT(dalpha_L3_j_3[1]), .SIGN_out(SIGN_dalpha_L3_j_3[1]));
SS_ADDSUB ADDSUB_dalpha_L3_1_4(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L3_j_4_netPar0[1], dalpha_L3_j_4_netPar1[1], dalpha_L3_j_4_netPar2[1] }), .SIGN({ SIGN_dalpha_L3_j_4_netPar0[1], SIGN_dalpha_L3_j_4_netPar1[1], SIGN_dalpha_L3_j_4_netPar2[1]}), .R_condition(rc[367]), .OUT(dalpha_L3_j_4[1]), .SIGN_out(SIGN_dalpha_L3_j_4[1]));
SS_ADDSUB ADDSUB_dalpha_L3_2_0(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L3_j_0_netPar0[2], dalpha_L3_j_0_netPar1[2], dalpha_L3_j_0_netPar2[2] }), .SIGN({ SIGN_dalpha_L3_j_0_netPar0[2], SIGN_dalpha_L3_j_0_netPar1[2], SIGN_dalpha_L3_j_0_netPar2[2]}), .R_condition(rc[368]), .OUT(dalpha_L3_j_0[2]), .SIGN_out(SIGN_dalpha_L3_j_0[2]));
SS_ADDSUB ADDSUB_dalpha_L3_2_1(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L3_j_1_netPar0[2], dalpha_L3_j_1_netPar1[2], dalpha_L3_j_1_netPar2[2] }), .SIGN({ SIGN_dalpha_L3_j_1_netPar0[2], SIGN_dalpha_L3_j_1_netPar1[2], SIGN_dalpha_L3_j_1_netPar2[2]}), .R_condition(rc[369]), .OUT(dalpha_L3_j_1[2]), .SIGN_out(SIGN_dalpha_L3_j_1[2]));
SS_ADDSUB ADDSUB_dalpha_L3_2_2(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L3_j_2_netPar0[2], dalpha_L3_j_2_netPar1[2], dalpha_L3_j_2_netPar2[2] }), .SIGN({ SIGN_dalpha_L3_j_2_netPar0[2], SIGN_dalpha_L3_j_2_netPar1[2], SIGN_dalpha_L3_j_2_netPar2[2]}), .R_condition(rc[370]), .OUT(dalpha_L3_j_2[2]), .SIGN_out(SIGN_dalpha_L3_j_2[2]));
SS_ADDSUB ADDSUB_dalpha_L3_2_3(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L3_j_3_netPar0[2], dalpha_L3_j_3_netPar1[2], dalpha_L3_j_3_netPar2[2] }), .SIGN({ SIGN_dalpha_L3_j_3_netPar0[2], SIGN_dalpha_L3_j_3_netPar1[2], SIGN_dalpha_L3_j_3_netPar2[2]}), .R_condition(rc[371]), .OUT(dalpha_L3_j_3[2]), .SIGN_out(SIGN_dalpha_L3_j_3[2]));
SS_ADDSUB ADDSUB_dalpha_L3_2_4(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L3_j_4_netPar0[2], dalpha_L3_j_4_netPar1[2], dalpha_L3_j_4_netPar2[2] }), .SIGN({ SIGN_dalpha_L3_j_4_netPar0[2], SIGN_dalpha_L3_j_4_netPar1[2], SIGN_dalpha_L3_j_4_netPar2[2]}), .R_condition(rc[372]), .OUT(dalpha_L3_j_4[2]), .SIGN_out(SIGN_dalpha_L3_j_4[2]));
SS_ADDSUB ADDSUB_dalpha_L3_3_0(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L3_j_0_netPar0[3], dalpha_L3_j_0_netPar1[3], dalpha_L3_j_0_netPar2[3] }), .SIGN({ SIGN_dalpha_L3_j_0_netPar0[3], SIGN_dalpha_L3_j_0_netPar1[3], SIGN_dalpha_L3_j_0_netPar2[3]}), .R_condition(rc[373]), .OUT(dalpha_L3_j_0[3]), .SIGN_out(SIGN_dalpha_L3_j_0[3]));
SS_ADDSUB ADDSUB_dalpha_L3_3_1(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L3_j_1_netPar0[3], dalpha_L3_j_1_netPar1[3], dalpha_L3_j_1_netPar2[3] }), .SIGN({ SIGN_dalpha_L3_j_1_netPar0[3], SIGN_dalpha_L3_j_1_netPar1[3], SIGN_dalpha_L3_j_1_netPar2[3]}), .R_condition(rc[374]), .OUT(dalpha_L3_j_1[3]), .SIGN_out(SIGN_dalpha_L3_j_1[3]));
SS_ADDSUB ADDSUB_dalpha_L3_3_2(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L3_j_2_netPar0[3], dalpha_L3_j_2_netPar1[3], dalpha_L3_j_2_netPar2[3] }), .SIGN({ SIGN_dalpha_L3_j_2_netPar0[3], SIGN_dalpha_L3_j_2_netPar1[3], SIGN_dalpha_L3_j_2_netPar2[3]}), .R_condition(rc[375]), .OUT(dalpha_L3_j_2[3]), .SIGN_out(SIGN_dalpha_L3_j_2[3]));
SS_ADDSUB ADDSUB_dalpha_L3_3_3(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L3_j_3_netPar0[3], dalpha_L3_j_3_netPar1[3], dalpha_L3_j_3_netPar2[3] }), .SIGN({ SIGN_dalpha_L3_j_3_netPar0[3], SIGN_dalpha_L3_j_3_netPar1[3], SIGN_dalpha_L3_j_3_netPar2[3]}), .R_condition(rc[376]), .OUT(dalpha_L3_j_3[3]), .SIGN_out(SIGN_dalpha_L3_j_3[3]));
SS_ADDSUB ADDSUB_dalpha_L3_3_4(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L3_j_4_netPar0[3], dalpha_L3_j_4_netPar1[3], dalpha_L3_j_4_netPar2[3] }), .SIGN({ SIGN_dalpha_L3_j_4_netPar0[3], SIGN_dalpha_L3_j_4_netPar1[3], SIGN_dalpha_L3_j_4_netPar2[3]}), .R_condition(rc[377]), .OUT(dalpha_L3_j_4[3]), .SIGN_out(SIGN_dalpha_L3_j_4[3]));
SS_ADDSUB ADDSUB_dalpha_L3_4_0(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L3_j_0_netPar0[4], dalpha_L3_j_0_netPar1[4], dalpha_L3_j_0_netPar2[4] }), .SIGN({ SIGN_dalpha_L3_j_0_netPar0[4], SIGN_dalpha_L3_j_0_netPar1[4], SIGN_dalpha_L3_j_0_netPar2[4]}), .R_condition(rc[378]), .OUT(dalpha_L3_j_0[4]), .SIGN_out(SIGN_dalpha_L3_j_0[4]));
SS_ADDSUB ADDSUB_dalpha_L3_4_1(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L3_j_1_netPar0[4], dalpha_L3_j_1_netPar1[4], dalpha_L3_j_1_netPar2[4] }), .SIGN({ SIGN_dalpha_L3_j_1_netPar0[4], SIGN_dalpha_L3_j_1_netPar1[4], SIGN_dalpha_L3_j_1_netPar2[4]}), .R_condition(rc[379]), .OUT(dalpha_L3_j_1[4]), .SIGN_out(SIGN_dalpha_L3_j_1[4]));
SS_ADDSUB ADDSUB_dalpha_L3_4_2(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L3_j_2_netPar0[4], dalpha_L3_j_2_netPar1[4], dalpha_L3_j_2_netPar2[4] }), .SIGN({ SIGN_dalpha_L3_j_2_netPar0[4], SIGN_dalpha_L3_j_2_netPar1[4], SIGN_dalpha_L3_j_2_netPar2[4]}), .R_condition(rc[380]), .OUT(dalpha_L3_j_2[4]), .SIGN_out(SIGN_dalpha_L3_j_2[4]));
SS_ADDSUB ADDSUB_dalpha_L3_4_3(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L3_j_3_netPar0[4], dalpha_L3_j_3_netPar1[4], dalpha_L3_j_3_netPar2[4] }), .SIGN({ SIGN_dalpha_L3_j_3_netPar0[4], SIGN_dalpha_L3_j_3_netPar1[4], SIGN_dalpha_L3_j_3_netPar2[4]}), .R_condition(rc[381]), .OUT(dalpha_L3_j_3[4]), .SIGN_out(SIGN_dalpha_L3_j_3[4]));
SS_ADDSUB ADDSUB_dalpha_L3_4_4(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L3_j_4_netPar0[4], dalpha_L3_j_4_netPar1[4], dalpha_L3_j_4_netPar2[4] }), .SIGN({ SIGN_dalpha_L3_j_4_netPar0[4], SIGN_dalpha_L3_j_4_netPar1[4], SIGN_dalpha_L3_j_4_netPar2[4]}), .R_condition(rc[382]), .OUT(dalpha_L3_j_4[4]), .SIGN_out(SIGN_dalpha_L3_j_4[4]));
SS_ADDSUB ADDSUB_dalpha_L3_5_0(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L3_j_0_netPar0[5], dalpha_L3_j_0_netPar1[5], dalpha_L3_j_0_netPar2[5] }), .SIGN({ SIGN_dalpha_L3_j_0_netPar0[5], SIGN_dalpha_L3_j_0_netPar1[5], SIGN_dalpha_L3_j_0_netPar2[5]}), .R_condition(rc[383]), .OUT(dalpha_L3_j_0[5]), .SIGN_out(SIGN_dalpha_L3_j_0[5]));
SS_ADDSUB ADDSUB_dalpha_L3_5_1(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L3_j_1_netPar0[5], dalpha_L3_j_1_netPar1[5], dalpha_L3_j_1_netPar2[5] }), .SIGN({ SIGN_dalpha_L3_j_1_netPar0[5], SIGN_dalpha_L3_j_1_netPar1[5], SIGN_dalpha_L3_j_1_netPar2[5]}), .R_condition(rc[384]), .OUT(dalpha_L3_j_1[5]), .SIGN_out(SIGN_dalpha_L3_j_1[5]));
SS_ADDSUB ADDSUB_dalpha_L3_5_2(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L3_j_2_netPar0[5], dalpha_L3_j_2_netPar1[5], dalpha_L3_j_2_netPar2[5] }), .SIGN({ SIGN_dalpha_L3_j_2_netPar0[5], SIGN_dalpha_L3_j_2_netPar1[5], SIGN_dalpha_L3_j_2_netPar2[5]}), .R_condition(rc[385]), .OUT(dalpha_L3_j_2[5]), .SIGN_out(SIGN_dalpha_L3_j_2[5]));
SS_ADDSUB ADDSUB_dalpha_L3_5_3(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L3_j_3_netPar0[5], dalpha_L3_j_3_netPar1[5], dalpha_L3_j_3_netPar2[5] }), .SIGN({ SIGN_dalpha_L3_j_3_netPar0[5], SIGN_dalpha_L3_j_3_netPar1[5], SIGN_dalpha_L3_j_3_netPar2[5]}), .R_condition(rc[386]), .OUT(dalpha_L3_j_3[5]), .SIGN_out(SIGN_dalpha_L3_j_3[5]));
SS_ADDSUB ADDSUB_dalpha_L3_5_4(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L3_j_4_netPar0[5], dalpha_L3_j_4_netPar1[5], dalpha_L3_j_4_netPar2[5] }), .SIGN({ SIGN_dalpha_L3_j_4_netPar0[5], SIGN_dalpha_L3_j_4_netPar1[5], SIGN_dalpha_L3_j_4_netPar2[5]}), .R_condition(rc[387]), .OUT(dalpha_L3_j_4[5]), .SIGN_out(SIGN_dalpha_L3_j_4[5]));
SS_ADDSUB ADDSUB_dalpha_L3_6_0(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L3_j_0_netPar0[6], dalpha_L3_j_0_netPar1[6], dalpha_L3_j_0_netPar2[6] }), .SIGN({ SIGN_dalpha_L3_j_0_netPar0[6], SIGN_dalpha_L3_j_0_netPar1[6], SIGN_dalpha_L3_j_0_netPar2[6]}), .R_condition(rc[388]), .OUT(dalpha_L3_j_0[6]), .SIGN_out(SIGN_dalpha_L3_j_0[6]));
SS_ADDSUB ADDSUB_dalpha_L3_6_1(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L3_j_1_netPar0[6], dalpha_L3_j_1_netPar1[6], dalpha_L3_j_1_netPar2[6] }), .SIGN({ SIGN_dalpha_L3_j_1_netPar0[6], SIGN_dalpha_L3_j_1_netPar1[6], SIGN_dalpha_L3_j_1_netPar2[6]}), .R_condition(rc[389]), .OUT(dalpha_L3_j_1[6]), .SIGN_out(SIGN_dalpha_L3_j_1[6]));
SS_ADDSUB ADDSUB_dalpha_L3_6_2(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L3_j_2_netPar0[6], dalpha_L3_j_2_netPar1[6], dalpha_L3_j_2_netPar2[6] }), .SIGN({ SIGN_dalpha_L3_j_2_netPar0[6], SIGN_dalpha_L3_j_2_netPar1[6], SIGN_dalpha_L3_j_2_netPar2[6]}), .R_condition(rc[390]), .OUT(dalpha_L3_j_2[6]), .SIGN_out(SIGN_dalpha_L3_j_2[6]));
SS_ADDSUB ADDSUB_dalpha_L3_6_3(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L3_j_3_netPar0[6], dalpha_L3_j_3_netPar1[6], dalpha_L3_j_3_netPar2[6] }), .SIGN({ SIGN_dalpha_L3_j_3_netPar0[6], SIGN_dalpha_L3_j_3_netPar1[6], SIGN_dalpha_L3_j_3_netPar2[6]}), .R_condition(rc[391]), .OUT(dalpha_L3_j_3[6]), .SIGN_out(SIGN_dalpha_L3_j_3[6]));
SS_ADDSUB ADDSUB_dalpha_L3_6_4(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L3_j_4_netPar0[6], dalpha_L3_j_4_netPar1[6], dalpha_L3_j_4_netPar2[6] }), .SIGN({ SIGN_dalpha_L3_j_4_netPar0[6], SIGN_dalpha_L3_j_4_netPar1[6], SIGN_dalpha_L3_j_4_netPar2[6]}), .R_condition(rc[392]), .OUT(dalpha_L3_j_4[6]), .SIGN_out(SIGN_dalpha_L3_j_4[6]));
SS_ADDSUB ADDSUB_dalpha_L3_7_0(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L3_j_0_netPar0[7], dalpha_L3_j_0_netPar1[7], dalpha_L3_j_0_netPar2[7] }), .SIGN({ SIGN_dalpha_L3_j_0_netPar0[7], SIGN_dalpha_L3_j_0_netPar1[7], SIGN_dalpha_L3_j_0_netPar2[7]}), .R_condition(rc[393]), .OUT(dalpha_L3_j_0[7]), .SIGN_out(SIGN_dalpha_L3_j_0[7]));
SS_ADDSUB ADDSUB_dalpha_L3_7_1(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L3_j_1_netPar0[7], dalpha_L3_j_1_netPar1[7], dalpha_L3_j_1_netPar2[7] }), .SIGN({ SIGN_dalpha_L3_j_1_netPar0[7], SIGN_dalpha_L3_j_1_netPar1[7], SIGN_dalpha_L3_j_1_netPar2[7]}), .R_condition(rc[394]), .OUT(dalpha_L3_j_1[7]), .SIGN_out(SIGN_dalpha_L3_j_1[7]));
SS_ADDSUB ADDSUB_dalpha_L3_7_2(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L3_j_2_netPar0[7], dalpha_L3_j_2_netPar1[7], dalpha_L3_j_2_netPar2[7] }), .SIGN({ SIGN_dalpha_L3_j_2_netPar0[7], SIGN_dalpha_L3_j_2_netPar1[7], SIGN_dalpha_L3_j_2_netPar2[7]}), .R_condition(rc[395]), .OUT(dalpha_L3_j_2[7]), .SIGN_out(SIGN_dalpha_L3_j_2[7]));
SS_ADDSUB ADDSUB_dalpha_L3_7_3(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L3_j_3_netPar0[7], dalpha_L3_j_3_netPar1[7], dalpha_L3_j_3_netPar2[7] }), .SIGN({ SIGN_dalpha_L3_j_3_netPar0[7], SIGN_dalpha_L3_j_3_netPar1[7], SIGN_dalpha_L3_j_3_netPar2[7]}), .R_condition(rc[396]), .OUT(dalpha_L3_j_3[7]), .SIGN_out(SIGN_dalpha_L3_j_3[7]));
SS_ADDSUB ADDSUB_dalpha_L3_7_4(.CLK(CLK), .INIT(INIT), .IN({ dalpha_L3_j_4_netPar0[7], dalpha_L3_j_4_netPar1[7], dalpha_L3_j_4_netPar2[7] }), .SIGN({ SIGN_dalpha_L3_j_4_netPar0[7], SIGN_dalpha_L3_j_4_netPar1[7], SIGN_dalpha_L3_j_4_netPar2[7]}), .R_condition(rc[397]), .OUT(dalpha_L3_j_4[7]), .SIGN_out(SIGN_dalpha_L3_j_4[7]));
defparam ADDSUB_dalpha_L3_0_0.N = 3;
defparam ADDSUB_dalpha_L3_0_1.N = 3;
defparam ADDSUB_dalpha_L3_0_2.N = 3;
defparam ADDSUB_dalpha_L3_0_3.N = 3;
defparam ADDSUB_dalpha_L3_0_4.N = 3;
defparam ADDSUB_dalpha_L3_1_0.N = 3;
defparam ADDSUB_dalpha_L3_1_1.N = 3;
defparam ADDSUB_dalpha_L3_1_2.N = 3;
defparam ADDSUB_dalpha_L3_1_3.N = 3;
defparam ADDSUB_dalpha_L3_1_4.N = 3;
defparam ADDSUB_dalpha_L3_2_0.N = 3;
defparam ADDSUB_dalpha_L3_2_1.N = 3;
defparam ADDSUB_dalpha_L3_2_2.N = 3;
defparam ADDSUB_dalpha_L3_2_3.N = 3;
defparam ADDSUB_dalpha_L3_2_4.N = 3;
defparam ADDSUB_dalpha_L3_3_0.N = 3;
defparam ADDSUB_dalpha_L3_3_1.N = 3;
defparam ADDSUB_dalpha_L3_3_2.N = 3;
defparam ADDSUB_dalpha_L3_3_3.N = 3;
defparam ADDSUB_dalpha_L3_3_4.N = 3;
defparam ADDSUB_dalpha_L3_4_0.N = 3;
defparam ADDSUB_dalpha_L3_4_1.N = 3;
defparam ADDSUB_dalpha_L3_4_2.N = 3;
defparam ADDSUB_dalpha_L3_4_3.N = 3;
defparam ADDSUB_dalpha_L3_4_4.N = 3;
defparam ADDSUB_dalpha_L3_5_0.N = 3;
defparam ADDSUB_dalpha_L3_5_1.N = 3;
defparam ADDSUB_dalpha_L3_5_2.N = 3;
defparam ADDSUB_dalpha_L3_5_3.N = 3;
defparam ADDSUB_dalpha_L3_5_4.N = 3;
defparam ADDSUB_dalpha_L3_6_0.N = 3;
defparam ADDSUB_dalpha_L3_6_1.N = 3;
defparam ADDSUB_dalpha_L3_6_2.N = 3;
defparam ADDSUB_dalpha_L3_6_3.N = 3;
defparam ADDSUB_dalpha_L3_6_4.N = 3;
defparam ADDSUB_dalpha_L3_7_0.N = 3;
defparam ADDSUB_dalpha_L3_7_1.N = 3;
defparam ADDSUB_dalpha_L3_7_2.N = 3;
defparam ADDSUB_dalpha_L3_7_3.N = 3;
defparam ADDSUB_dalpha_L3_7_4.N = 3;
defparam ADDSUB_dalpha_L3_0_0.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L3_0_1.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L3_0_2.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L3_0_3.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L3_0_4.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L3_1_0.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L3_1_1.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L3_1_2.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L3_1_3.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L3_1_4.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L3_2_0.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L3_2_1.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L3_2_2.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L3_2_3.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L3_2_4.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L3_3_0.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L3_3_1.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L3_3_2.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L3_3_3.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L3_3_4.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L3_4_0.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L3_4_1.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L3_4_2.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L3_4_3.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L3_4_4.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L3_5_0.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L3_5_1.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L3_5_2.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L3_5_3.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L3_5_4.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L3_6_0.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L3_6_1.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L3_6_2.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L3_6_3.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L3_6_4.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L3_7_0.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L3_7_1.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L3_7_2.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L3_7_3.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dalpha_L3_7_4.DIFFCOUNTER_SIZE = 3;

SS_ADDSUB ADDSUB_dbeta_L3_0(.CLK(CLK), .INIT(INIT), .IN({ dbeta_L3_netPar0[0], dbeta_L3_netPar1[0], dbeta_L3_netPar2[0] }), .SIGN({ SIGN_dbeta_L3_netPar0[0], SIGN_dbeta_L3_netPar1[0], SIGN_dbeta_L3_netPar2[0]}), .R_condition(rc[398]), .OUT(dbeta_L3[0]), .SIGN_out(SIGN_dbeta_L3[0]));
SS_ADDSUB ADDSUB_dbeta_L3_1(.CLK(CLK), .INIT(INIT), .IN({ dbeta_L3_netPar0[1], dbeta_L3_netPar1[1], dbeta_L3_netPar2[1] }), .SIGN({ SIGN_dbeta_L3_netPar0[1], SIGN_dbeta_L3_netPar1[1], SIGN_dbeta_L3_netPar2[1]}), .R_condition(rc[399]), .OUT(dbeta_L3[1]), .SIGN_out(SIGN_dbeta_L3[1]));
SS_ADDSUB ADDSUB_dbeta_L3_2(.CLK(CLK), .INIT(INIT), .IN({ dbeta_L3_netPar0[2], dbeta_L3_netPar1[2], dbeta_L3_netPar2[2] }), .SIGN({ SIGN_dbeta_L3_netPar0[2], SIGN_dbeta_L3_netPar1[2], SIGN_dbeta_L3_netPar2[2]}), .R_condition(rc[400]), .OUT(dbeta_L3[2]), .SIGN_out(SIGN_dbeta_L3[2]));
SS_ADDSUB ADDSUB_dbeta_L3_3(.CLK(CLK), .INIT(INIT), .IN({ dbeta_L3_netPar0[3], dbeta_L3_netPar1[3], dbeta_L3_netPar2[3] }), .SIGN({ SIGN_dbeta_L3_netPar0[3], SIGN_dbeta_L3_netPar1[3], SIGN_dbeta_L3_netPar2[3]}), .R_condition(rc[401]), .OUT(dbeta_L3[3]), .SIGN_out(SIGN_dbeta_L3[3]));
SS_ADDSUB ADDSUB_dbeta_L3_4(.CLK(CLK), .INIT(INIT), .IN({ dbeta_L3_netPar0[4], dbeta_L3_netPar1[4], dbeta_L3_netPar2[4] }), .SIGN({ SIGN_dbeta_L3_netPar0[4], SIGN_dbeta_L3_netPar1[4], SIGN_dbeta_L3_netPar2[4]}), .R_condition(rc[402]), .OUT(dbeta_L3[4]), .SIGN_out(SIGN_dbeta_L3[4]));
defparam ADDSUB_dbeta_L3_0.N = 3;
defparam ADDSUB_dbeta_L3_1.N = 3;
defparam ADDSUB_dbeta_L3_2.N = 3;
defparam ADDSUB_dbeta_L3_3.N = 3;
defparam ADDSUB_dbeta_L3_4.N = 3;
defparam ADDSUB_dbeta_L3_0.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dbeta_L3_1.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dbeta_L3_2.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dbeta_L3_3.DIFFCOUNTER_SIZE = 3;
defparam ADDSUB_dbeta_L3_4.DIFFCOUNTER_SIZE = 3;



endmodule
