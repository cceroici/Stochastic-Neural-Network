// Chris Ceroici

// LFSR seed signals for 16 bit LFSRs

module SEED(INIT,S0,S2,S4,S6,S8,S10,S12,S14,S16,S18,S20,S22,S24,S26,S28,S30,S32,S34,S36,S38,S40,S42,S44,S46,S48,S50,S52,S54,S56,S58,S60,S62,S64,S66,S68,S70,S72,S74,S76,S78,S80,S82,S84,S86,S88,S90,S92,S94,S96,S98,S100,S102,S104,S106,S108,S110,S112,S114,S116,S118,S120,S122,S124,S126,S128,S130,S132,S134,S136,S138,S140,S142,S144,S146,S148,S150,S152,S154,S156,S158,S160,S162,S164,S166,S168,S170,S172,S174,S176,S178,S180,S182,S184,S186,S188,S190,S192,S194,S196,S198,S200,S202,S204,S206,S208,S210,S212,S214,S216,S218,S220,S222,S224,S226,S228,S230,S232,S234,S236,S238,S240,S242,S244,S246,S248,S250,S252,S254,S256,S258,S260,S262,S264,S266,S268,S270,S272,S274,S276,S278,S1,S3,S5,S7,S9,S11,S13,S15,S17,S19,S21,S23,S25,S27,S29,S31,S33,S35,S37,S39,S41,S43,S45,S47,S49,S51,S53,S55,S57,S59,S61,S63,S65,S67,S69,S71,S73,S75,S77,S79,S81,S83,S85,S87,S89,S91,S93,S95,S97,S99,S101,S103,S105,S107,S109,S111,S113,S115,S117,S119,S121,S123,S125,S127,S129,S131,S133,S135,S137,S139,S141,S143,S145,S147,S149,S151,S153,S155,S157,S159,S161,S163,S165,S167,S169,S171,S173,S175,S177,S179,S181,S183,S185,S187,S189,S191,S193,S195,S197,S199,S201,S203,S205,S207,S209,S211,S213,S215,S217,S219,S221,S223,S225,S227,S229,S231,S233,S235,S237,S239,S241,S243,S245,S247,S249,S251,S253,S255,S257,S259,S261,S263,S265,S267,S269,S271,S273,S275,S277,S279);

parameter LFSR_S = 16; // LFSR size

input INIT; // Initialization signal (new set)

output [LFSR_S-1:0] S0,S1,S2,S3,S4,S5,S6,S7,S8,S9,S10,S11,S12,S13,S14,S15,S16,S17,S18,S19,S20,S21,S22,S23,S24,S25,S26,S27,S28,S29,S30,S31,S32,S33,S34,S35,S36,S37,S38,S39,S40,S41,S42,S43,S44,S45,S46,S47,S48,S49,S50,S51,S52,S53,S54,S55,S56,S57,S58,S59,S60,S61,S62,S63,S64,S65,S66,S67,S68,S69,S70,S71,S72,S73,S74,S75,S76,S77,S78,S79,S80,S81,S82,S83,S84,S85,S86,S87,S88,S89,S90,S91,S92,S93,S94,S95,S96,S97,S98,S99,S100,S101,S102,S103,S104,S105,S106,S107,S108,S109,S110,S111,S112,S113,S114,S115,S116,S117,S118,S119,S120,S121,S122,S123,S124,S125,S126,S127,S128,S129,S130,S131,S132,S133,S134,S135,S136,S137,S138,S139,S140,S141,S142,S143,S144,S145,S146,S147,S148,S149,S150,S151,S152,S153,S154,S155,S156,S157,S158,S159,S160,S161,S162,S163,S164,S165,S166,S167,S168,S169,S170,S171,S172,S173,S174,S175,S176,S177,S178,S179,S180,S181,S182,S183,S184,S185,S186,S187,S188,S189,S190,S191,S192,S193,S194,S195,S196,S197,S198,S199,S200,S201,S202,S203,S204,S205,S206,S207,S208,S209,S210,S211,S212,S213,S214,S215,S216,S217,S218,S219,S220,S221,S222,S223,S224,S225,S226,S227,S228,S229,S230,S231,S232,S233,S234,S235,S236,S237,S238,S239,S240,S241,S242,S243,S244,S245,S246,S247,S248,S249,S250,S251,S252,S253,S254,S255,S256,S257,S258,S259,S260,S261,S262,S263,S264,S265,S266,S267,S268,S269,S270,S271,S272,S273,S274,S275,S276,S277,S278,S279;

integer n1 = 0; // Set counter (Decoder)
integer n2 = 0; // Set counter (Channel simulator)
integer ndiff = 1; // differential counter

// Set 1 Seeds: 
reg [LFSR_S-1:0] S0reg = 16'b0001000001011000;
reg [LFSR_S-1:0] S1reg = 16'b0011111110011011;
reg [LFSR_S-1:0] S2reg = 16'b1011010010000000;
reg [LFSR_S-1:0] S3reg = 16'b0110110011010010;
reg [LFSR_S-1:0] S4reg = 16'b1011101010010100;
reg [LFSR_S-1:0] S5reg = 16'b1101010101100110;
reg [LFSR_S-1:0] S6reg = 16'b1101100101011010;
reg [LFSR_S-1:0] S7reg = 16'b1110111011011011;
reg [LFSR_S-1:0] S8reg = 16'b0011110010011100;
reg [LFSR_S-1:0] S9reg = 16'b1001010000001000;
reg [LFSR_S-1:0] S10reg = 16'b1111101101000011;
reg [LFSR_S-1:0] S11reg = 16'b1100101100100001;
reg [LFSR_S-1:0] S12reg = 16'b0011000100011100;
reg [LFSR_S-1:0] S13reg = 16'b1010000000000010;
reg [LFSR_S-1:0] S14reg = 16'b0100111101100011;
reg [LFSR_S-1:0] S15reg = 16'b1001010101100111;
reg [LFSR_S-1:0] S16reg = 16'b1000000101100000;
reg [LFSR_S-1:0] S17reg = 16'b0110000100111110;
reg [LFSR_S-1:0] S18reg = 16'b1000010100110011;
reg [LFSR_S-1:0] S19reg = 16'b0101101010000001;
reg [LFSR_S-1:0] S20reg = 16'b1111011100001001;
reg [LFSR_S-1:0] S21reg = 16'b0110011100101011;
reg [LFSR_S-1:0] S22reg = 16'b0100110110011000;
reg [LFSR_S-1:0] S23reg = 16'b1011111011101101;
reg [LFSR_S-1:0] S24reg = 16'b0010101100111111;
reg [LFSR_S-1:0] S25reg = 16'b1101010001001110;
reg [LFSR_S-1:0] S26reg = 16'b1100111000100101;
reg [LFSR_S-1:0] S27reg = 16'b1001111000100101;
reg [LFSR_S-1:0] S28reg = 16'b0011110111010110;
reg [LFSR_S-1:0] S29reg = 16'b0010000111110101;
reg [LFSR_S-1:0] S30reg = 16'b0110100001100101;
reg [LFSR_S-1:0] S31reg = 16'b1010100100100100;
reg [LFSR_S-1:0] S32reg = 16'b1111001100101000;
reg [LFSR_S-1:0] S33reg = 16'b1111010000111111;
reg [LFSR_S-1:0] S34reg = 16'b1001011110110010;
reg [LFSR_S-1:0] S35reg = 16'b0101110110000001;
reg [LFSR_S-1:0] S36reg = 16'b0101010001001101;
reg [LFSR_S-1:0] S37reg = 16'b1000010101001000;
reg [LFSR_S-1:0] S38reg = 16'b0111111101000100;
reg [LFSR_S-1:0] S39reg = 16'b1110110110101101;
reg [LFSR_S-1:0] S40reg = 16'b1010001101100111;
reg [LFSR_S-1:0] S41reg = 16'b0110011100011100;
reg [LFSR_S-1:0] S42reg = 16'b1011000011101000;
reg [LFSR_S-1:0] S43reg = 16'b1110011001000111;
reg [LFSR_S-1:0] S44reg = 16'b1000000010000110;
reg [LFSR_S-1:0] S45reg = 16'b1110010011000010;
reg [LFSR_S-1:0] S46reg = 16'b1101111110111101;
reg [LFSR_S-1:0] S47reg = 16'b0100100010100110;
reg [LFSR_S-1:0] S48reg = 16'b1101110001101110;
reg [LFSR_S-1:0] S49reg = 16'b1101110111100101;
reg [LFSR_S-1:0] S50reg = 16'b0010001010010111;
reg [LFSR_S-1:0] S51reg = 16'b1101001000111111;
reg [LFSR_S-1:0] S52reg = 16'b0000000001001000;
reg [LFSR_S-1:0] S53reg = 16'b1110011011110101;
reg [LFSR_S-1:0] S54reg = 16'b1111001010011000;
reg [LFSR_S-1:0] S55reg = 16'b0101100110000100;
reg [LFSR_S-1:0] S56reg = 16'b1010111010111111;
reg [LFSR_S-1:0] S57reg = 16'b1100000110011001;
reg [LFSR_S-1:0] S58reg = 16'b0011101010001010;
reg [LFSR_S-1:0] S59reg = 16'b1001111100000111;
reg [LFSR_S-1:0] S60reg = 16'b1111100111000010;
reg [LFSR_S-1:0] S61reg = 16'b1010011101100000;
reg [LFSR_S-1:0] S62reg = 16'b0000001000001100;
reg [LFSR_S-1:0] S63reg = 16'b1110111110100001;
reg [LFSR_S-1:0] S64reg = 16'b1111111111101001;
reg [LFSR_S-1:0] S65reg = 16'b1011110001100010;
reg [LFSR_S-1:0] S66reg = 16'b1110000111110011;
reg [LFSR_S-1:0] S67reg = 16'b1000011011100101;
reg [LFSR_S-1:0] S68reg = 16'b0101111101100010;
reg [LFSR_S-1:0] S69reg = 16'b0010001001001000;
reg [LFSR_S-1:0] S70reg = 16'b0011111001000111;
reg [LFSR_S-1:0] S71reg = 16'b1011000111001000;
reg [LFSR_S-1:0] S72reg = 16'b1111000010111101;
reg [LFSR_S-1:0] S73reg = 16'b0111001101111111;
reg [LFSR_S-1:0] S74reg = 16'b0110110001100000;
reg [LFSR_S-1:0] S75reg = 16'b0110111000110000;
reg [LFSR_S-1:0] S76reg = 16'b1100110101110001;
reg [LFSR_S-1:0] S77reg = 16'b1011010001010101;
reg [LFSR_S-1:0] S78reg = 16'b0110001001101111;
reg [LFSR_S-1:0] S79reg = 16'b0001010000010110;
reg [LFSR_S-1:0] S80reg = 16'b1110010111000111;
reg [LFSR_S-1:0] S81reg = 16'b0101110010100010;
reg [LFSR_S-1:0] S82reg = 16'b0110001011110000;
reg [LFSR_S-1:0] S83reg = 16'b1100000010000011;
reg [LFSR_S-1:0] S84reg = 16'b1001001101101111;
reg [LFSR_S-1:0] S85reg = 16'b1011011101101101;
reg [LFSR_S-1:0] S86reg = 16'b1010001100110001;
reg [LFSR_S-1:0] S87reg = 16'b1000011000110011;
reg [LFSR_S-1:0] S88reg = 16'b0001000011101000;
reg [LFSR_S-1:0] S89reg = 16'b1110110010011111;
reg [LFSR_S-1:0] S90reg = 16'b1100011111100101;
reg [LFSR_S-1:0] S91reg = 16'b1100001101010111;
reg [LFSR_S-1:0] S92reg = 16'b0001010101000001;
reg [LFSR_S-1:0] S93reg = 16'b1101010111111100;
reg [LFSR_S-1:0] S94reg = 16'b1100011011000100;
reg [LFSR_S-1:0] S95reg = 16'b0101001100010010;
reg [LFSR_S-1:0] S96reg = 16'b1111100101010011;
reg [LFSR_S-1:0] S97reg = 16'b1100110011011111;
reg [LFSR_S-1:0] S98reg = 16'b0110001101000000;
reg [LFSR_S-1:0] S99reg = 16'b1000111000011001;
reg [LFSR_S-1:0] S100reg = 16'b1111101111011111;
reg [LFSR_S-1:0] S101reg = 16'b1101011000011001;
reg [LFSR_S-1:0] S102reg = 16'b1010011111101010;
reg [LFSR_S-1:0] S103reg = 16'b0111010111001111;
reg [LFSR_S-1:0] S104reg = 16'b0100011001111000;
reg [LFSR_S-1:0] S105reg = 16'b0100011111100010;
reg [LFSR_S-1:0] S106reg = 16'b0011101010100010;
reg [LFSR_S-1:0] S107reg = 16'b1011010001100100;
reg [LFSR_S-1:0] S108reg = 16'b1101001110001001;
reg [LFSR_S-1:0] S109reg = 16'b1011100001110101;
reg [LFSR_S-1:0] S110reg = 16'b0101000011110101;
reg [LFSR_S-1:0] S111reg = 16'b0011110001110100;
reg [LFSR_S-1:0] S112reg = 16'b0001001100011110;
reg [LFSR_S-1:0] S113reg = 16'b1010010110011101;
reg [LFSR_S-1:0] S114reg = 16'b1111001110110111;
reg [LFSR_S-1:0] S115reg = 16'b0110011110010000;
reg [LFSR_S-1:0] S116reg = 16'b1110111111100000;
reg [LFSR_S-1:0] S117reg = 16'b1100101111001011;
reg [LFSR_S-1:0] S118reg = 16'b0000000001100100;
reg [LFSR_S-1:0] S119reg = 16'b0010000010111111;
reg [LFSR_S-1:0] S120reg = 16'b1100100101000011;
reg [LFSR_S-1:0] S121reg = 16'b1010000111000001;
reg [LFSR_S-1:0] S122reg = 16'b1100111011010011;
reg [LFSR_S-1:0] S123reg = 16'b1100010011010101;
reg [LFSR_S-1:0] S124reg = 16'b1101110001000101;
reg [LFSR_S-1:0] S125reg = 16'b0110011001000110;
reg [LFSR_S-1:0] S126reg = 16'b1100100000110101;
reg [LFSR_S-1:0] S127reg = 16'b1001000001110110;
reg [LFSR_S-1:0] S128reg = 16'b1100101011100101;
reg [LFSR_S-1:0] S129reg = 16'b1011000100010010;
reg [LFSR_S-1:0] S130reg = 16'b1011111001110100;
reg [LFSR_S-1:0] S131reg = 16'b1010001000000000;
reg [LFSR_S-1:0] S132reg = 16'b1010111000100010;
reg [LFSR_S-1:0] S133reg = 16'b0010010001111010;
reg [LFSR_S-1:0] S134reg = 16'b1011011100110100;
reg [LFSR_S-1:0] S135reg = 16'b1010010101001100;
reg [LFSR_S-1:0] S136reg = 16'b0111000101000101;
reg [LFSR_S-1:0] S137reg = 16'b1111001111001101;
reg [LFSR_S-1:0] S138reg = 16'b0110011010010000;
reg [LFSR_S-1:0] S139reg = 16'b1101100101011001;
reg [LFSR_S-1:0] S140reg = 16'b0010000100101001;
reg [LFSR_S-1:0] S141reg = 16'b0111101100101101;
reg [LFSR_S-1:0] S142reg = 16'b1010111101101101;
reg [LFSR_S-1:0] S143reg = 16'b0001100101010010;
reg [LFSR_S-1:0] S144reg = 16'b1100110010110001;
reg [LFSR_S-1:0] S145reg = 16'b0110100000111000;
reg [LFSR_S-1:0] S146reg = 16'b1100000010100101;
reg [LFSR_S-1:0] S147reg = 16'b1001100011110101;
reg [LFSR_S-1:0] S148reg = 16'b1100000011110101;
reg [LFSR_S-1:0] S149reg = 16'b1000111100111001;
reg [LFSR_S-1:0] S150reg = 16'b1111011001011100;
reg [LFSR_S-1:0] S151reg = 16'b1110100110100111;
reg [LFSR_S-1:0] S152reg = 16'b1001101100001011;
reg [LFSR_S-1:0] S153reg = 16'b0010101011100010;
reg [LFSR_S-1:0] S154reg = 16'b1111010010101001;
reg [LFSR_S-1:0] S155reg = 16'b0100010100001111;
reg [LFSR_S-1:0] S156reg = 16'b0110110001101110;
reg [LFSR_S-1:0] S157reg = 16'b0000011101110111;
reg [LFSR_S-1:0] S158reg = 16'b1001100101110010;
reg [LFSR_S-1:0] S159reg = 16'b1011011001010000;
reg [LFSR_S-1:0] S160reg = 16'b1100000011000001;
reg [LFSR_S-1:0] S161reg = 16'b1101011011111001;
reg [LFSR_S-1:0] S162reg = 16'b0101101101001110;
reg [LFSR_S-1:0] S163reg = 16'b0001010100101010;
reg [LFSR_S-1:0] S164reg = 16'b1101000100100100;
reg [LFSR_S-1:0] S165reg = 16'b0100000011001001;
reg [LFSR_S-1:0] S166reg = 16'b0001110101110010;
reg [LFSR_S-1:0] S167reg = 16'b1101010011101011;
reg [LFSR_S-1:0] S168reg = 16'b1011100100110101;
reg [LFSR_S-1:0] S169reg = 16'b0111100010010100;
reg [LFSR_S-1:0] S170reg = 16'b1010001011001011;
reg [LFSR_S-1:0] S171reg = 16'b1101010101100011;
reg [LFSR_S-1:0] S172reg = 16'b1110000011000010;
reg [LFSR_S-1:0] S173reg = 16'b0111001111100001;
reg [LFSR_S-1:0] S174reg = 16'b1000000011000111;
reg [LFSR_S-1:0] S175reg = 16'b0110101011111010;
reg [LFSR_S-1:0] S176reg = 16'b1011101011001111;
reg [LFSR_S-1:0] S177reg = 16'b1111000110000000;
reg [LFSR_S-1:0] S178reg = 16'b1100001111001100;
reg [LFSR_S-1:0] S179reg = 16'b0010101000011101;
reg [LFSR_S-1:0] S180reg = 16'b1000101010001101;
reg [LFSR_S-1:0] S181reg = 16'b1101100001111000;
reg [LFSR_S-1:0] S182reg = 16'b0000011100111101;
reg [LFSR_S-1:0] S183reg = 16'b0101001111011101;
reg [LFSR_S-1:0] S184reg = 16'b0011100011100000;
reg [LFSR_S-1:0] S185reg = 16'b0110000001000110;
reg [LFSR_S-1:0] S186reg = 16'b0111111011100111;
reg [LFSR_S-1:0] S187reg = 16'b1010010011110010;
reg [LFSR_S-1:0] S188reg = 16'b1010000110011011;
reg [LFSR_S-1:0] S189reg = 16'b0010011100111111;
reg [LFSR_S-1:0] S190reg = 16'b0010000001011101;
reg [LFSR_S-1:0] S191reg = 16'b0000111000111000;
reg [LFSR_S-1:0] S192reg = 16'b1110010010011110;
reg [LFSR_S-1:0] S193reg = 16'b0100101011111100;
reg [LFSR_S-1:0] S194reg = 16'b0101011001111100;
reg [LFSR_S-1:0] S195reg = 16'b0110011001011010;
reg [LFSR_S-1:0] S196reg = 16'b1000111111001111;
reg [LFSR_S-1:0] S197reg = 16'b0011100111110100;
reg [LFSR_S-1:0] S198reg = 16'b1101010100100011;
reg [LFSR_S-1:0] S199reg = 16'b1110000101011101;
reg [LFSR_S-1:0] S200reg = 16'b1101111100011101;
reg [LFSR_S-1:0] S201reg = 16'b0000101100001000;
reg [LFSR_S-1:0] S202reg = 16'b0110001001111101;
reg [LFSR_S-1:0] S203reg = 16'b1110000000100100;
reg [LFSR_S-1:0] S204reg = 16'b0100000101010100;
reg [LFSR_S-1:0] S205reg = 16'b0110001011011010;
reg [LFSR_S-1:0] S206reg = 16'b1101000111100101;
reg [LFSR_S-1:0] S207reg = 16'b1010111001011111;
reg [LFSR_S-1:0] S208reg = 16'b0010101100010110;
reg [LFSR_S-1:0] S209reg = 16'b1101101101000101;
reg [LFSR_S-1:0] S210reg = 16'b0110001100001110;
reg [LFSR_S-1:0] S211reg = 16'b0000010111011001;
reg [LFSR_S-1:0] S212reg = 16'b0010110100011110;
reg [LFSR_S-1:0] S213reg = 16'b0010100100000111;
reg [LFSR_S-1:0] S214reg = 16'b0001001111011010;
reg [LFSR_S-1:0] S215reg = 16'b1001111111111111;
reg [LFSR_S-1:0] S216reg = 16'b1100010000000000;
reg [LFSR_S-1:0] S217reg = 16'b0110001001001100;
reg [LFSR_S-1:0] S218reg = 16'b0011001001111000;
reg [LFSR_S-1:0] S219reg = 16'b0111101111100101;
reg [LFSR_S-1:0] S220reg = 16'b0101110010011110;
reg [LFSR_S-1:0] S221reg = 16'b1101110110111001;
reg [LFSR_S-1:0] S222reg = 16'b0011100100110111;
reg [LFSR_S-1:0] S223reg = 16'b1001001010111111;
reg [LFSR_S-1:0] S224reg = 16'b1010011001100111;
reg [LFSR_S-1:0] S225reg = 16'b0000011111100010;
reg [LFSR_S-1:0] S226reg = 16'b0111100001011111;
reg [LFSR_S-1:0] S227reg = 16'b1011101000010000;
reg [LFSR_S-1:0] S228reg = 16'b0111101000111010;
reg [LFSR_S-1:0] S229reg = 16'b1001101101110011;
reg [LFSR_S-1:0] S230reg = 16'b0110000010111000;
reg [LFSR_S-1:0] S231reg = 16'b1010110001010101;
reg [LFSR_S-1:0] S232reg = 16'b1101011111000001;
reg [LFSR_S-1:0] S233reg = 16'b0000101011000010;
reg [LFSR_S-1:0] S234reg = 16'b1011100000100110;
reg [LFSR_S-1:0] S235reg = 16'b1001001010000001;
reg [LFSR_S-1:0] S236reg = 16'b0111010111001000;
reg [LFSR_S-1:0] S237reg = 16'b1111110101011000;
reg [LFSR_S-1:0] S238reg = 16'b1001001000000011;
reg [LFSR_S-1:0] S239reg = 16'b1101000101000011;
reg [LFSR_S-1:0] S240reg = 16'b1111000100011110;
reg [LFSR_S-1:0] S241reg = 16'b0001010111010000;
reg [LFSR_S-1:0] S242reg = 16'b0010111001010000;
reg [LFSR_S-1:0] S243reg = 16'b0010011001010000;
reg [LFSR_S-1:0] S244reg = 16'b1000110010111110;
reg [LFSR_S-1:0] S245reg = 16'b1010110111000000;
reg [LFSR_S-1:0] S246reg = 16'b1101010000011101;
reg [LFSR_S-1:0] S247reg = 16'b1000101100110010;
reg [LFSR_S-1:0] S248reg = 16'b1101010101010011;
reg [LFSR_S-1:0] S249reg = 16'b0100011011100000;
reg [LFSR_S-1:0] S250reg = 16'b1011001010101101;
reg [LFSR_S-1:0] S251reg = 16'b1110000101100111;
reg [LFSR_S-1:0] S252reg = 16'b0010010010111010;
reg [LFSR_S-1:0] S253reg = 16'b0111101101110000;
reg [LFSR_S-1:0] S254reg = 16'b0101001011010001;
reg [LFSR_S-1:0] S255reg = 16'b1010110001100100;
reg [LFSR_S-1:0] S256reg = 16'b0111010011000110;
reg [LFSR_S-1:0] S257reg = 16'b0010010110001110;
reg [LFSR_S-1:0] S258reg = 16'b1001010001000001;
reg [LFSR_S-1:0] S259reg = 16'b0110001000011000;
reg [LFSR_S-1:0] S260reg = 16'b1011011100001000;
reg [LFSR_S-1:0] S261reg = 16'b1100100011011000;
reg [LFSR_S-1:0] S262reg = 16'b0101001001101110;
reg [LFSR_S-1:0] S263reg = 16'b1110000101100000;
reg [LFSR_S-1:0] S264reg = 16'b0100010100001010;
reg [LFSR_S-1:0] S265reg = 16'b0001100001010111;
reg [LFSR_S-1:0] S266reg = 16'b0111111000110001;
reg [LFSR_S-1:0] S267reg = 16'b0011100001101010;
reg [LFSR_S-1:0] S268reg = 16'b1100100010100101;
reg [LFSR_S-1:0] S269reg = 16'b1100100110000010;
reg [LFSR_S-1:0] S270reg = 16'b1000100010100111;
reg [LFSR_S-1:0] S271reg = 16'b1101110000010111;
reg [LFSR_S-1:0] S272reg = 16'b0110101101110010;
reg [LFSR_S-1:0] S273reg = 16'b0110100000001000;
reg [LFSR_S-1:0] S274reg = 16'b0011011010100000;
reg [LFSR_S-1:0] S275reg = 16'b1110101100101111;
reg [LFSR_S-1:0] S276reg = 16'b1001000000101100;
reg [LFSR_S-1:0] S277reg = 16'b0111010000010110;
reg [LFSR_S-1:0] S278reg = 16'b0000001000101010;
reg [LFSR_S-1:0] S279reg = 16'b1111010111001011;

assign S0[LFSR_S-1:0] = S0reg;
assign S1[LFSR_S-1:0] = S1reg;
assign S2[LFSR_S-1:0] = S2reg;
assign S3[LFSR_S-1:0] = S3reg;
assign S4[LFSR_S-1:0] = S4reg;
assign S5[LFSR_S-1:0] = S5reg;
assign S6[LFSR_S-1:0] = S6reg;
assign S7[LFSR_S-1:0] = S7reg;
assign S8[LFSR_S-1:0] = S8reg;
assign S9[LFSR_S-1:0] = S9reg;
assign S10[LFSR_S-1:0] = S10reg;
assign S11[LFSR_S-1:0] = S11reg;
assign S12[LFSR_S-1:0] = S12reg;
assign S13[LFSR_S-1:0] = S13reg;
assign S14[LFSR_S-1:0] = S14reg;
assign S15[LFSR_S-1:0] = S15reg;
assign S16[LFSR_S-1:0] = S16reg;
assign S17[LFSR_S-1:0] = S17reg;
assign S18[LFSR_S-1:0] = S18reg;
assign S19[LFSR_S-1:0] = S19reg;
assign S20[LFSR_S-1:0] = S20reg;
assign S21[LFSR_S-1:0] = S21reg;
assign S22[LFSR_S-1:0] = S22reg;
assign S23[LFSR_S-1:0] = S23reg;
assign S24[LFSR_S-1:0] = S24reg;
assign S25[LFSR_S-1:0] = S25reg;
assign S26[LFSR_S-1:0] = S26reg;
assign S27[LFSR_S-1:0] = S27reg;
assign S28[LFSR_S-1:0] = S28reg;
assign S29[LFSR_S-1:0] = S29reg;
assign S30[LFSR_S-1:0] = S30reg;
assign S31[LFSR_S-1:0] = S31reg;
assign S32[LFSR_S-1:0] = S32reg;
assign S33[LFSR_S-1:0] = S33reg;
assign S34[LFSR_S-1:0] = S34reg;
assign S35[LFSR_S-1:0] = S35reg;
assign S36[LFSR_S-1:0] = S36reg;
assign S37[LFSR_S-1:0] = S37reg;
assign S38[LFSR_S-1:0] = S38reg;
assign S39[LFSR_S-1:0] = S39reg;
assign S40[LFSR_S-1:0] = S40reg;
assign S41[LFSR_S-1:0] = S41reg;
assign S42[LFSR_S-1:0] = S42reg;
assign S43[LFSR_S-1:0] = S43reg;
assign S44[LFSR_S-1:0] = S44reg;
assign S45[LFSR_S-1:0] = S45reg;
assign S46[LFSR_S-1:0] = S46reg;
assign S47[LFSR_S-1:0] = S47reg;
assign S48[LFSR_S-1:0] = S48reg;
assign S49[LFSR_S-1:0] = S49reg;
assign S50[LFSR_S-1:0] = S50reg;
assign S51[LFSR_S-1:0] = S51reg;
assign S52[LFSR_S-1:0] = S52reg;
assign S53[LFSR_S-1:0] = S53reg;
assign S54[LFSR_S-1:0] = S54reg;
assign S55[LFSR_S-1:0] = S55reg;
assign S56[LFSR_S-1:0] = S56reg;
assign S57[LFSR_S-1:0] = S57reg;
assign S58[LFSR_S-1:0] = S58reg;
assign S59[LFSR_S-1:0] = S59reg;
assign S60[LFSR_S-1:0] = S60reg;
assign S61[LFSR_S-1:0] = S61reg;
assign S62[LFSR_S-1:0] = S62reg;
assign S63[LFSR_S-1:0] = S63reg;
assign S64[LFSR_S-1:0] = S64reg;
assign S65[LFSR_S-1:0] = S65reg;
assign S66[LFSR_S-1:0] = S66reg;
assign S67[LFSR_S-1:0] = S67reg;
assign S68[LFSR_S-1:0] = S68reg;
assign S69[LFSR_S-1:0] = S69reg;
assign S70[LFSR_S-1:0] = S70reg;
assign S71[LFSR_S-1:0] = S71reg;
assign S72[LFSR_S-1:0] = S72reg;
assign S73[LFSR_S-1:0] = S73reg;
assign S74[LFSR_S-1:0] = S74reg;
assign S75[LFSR_S-1:0] = S75reg;
assign S76[LFSR_S-1:0] = S76reg;
assign S77[LFSR_S-1:0] = S77reg;
assign S78[LFSR_S-1:0] = S78reg;
assign S79[LFSR_S-1:0] = S79reg;
assign S80[LFSR_S-1:0] = S80reg;
assign S81[LFSR_S-1:0] = S81reg;
assign S82[LFSR_S-1:0] = S82reg;
assign S83[LFSR_S-1:0] = S83reg;
assign S84[LFSR_S-1:0] = S84reg;
assign S85[LFSR_S-1:0] = S85reg;
assign S86[LFSR_S-1:0] = S86reg;
assign S87[LFSR_S-1:0] = S87reg;
assign S88[LFSR_S-1:0] = S88reg;
assign S89[LFSR_S-1:0] = S89reg;
assign S90[LFSR_S-1:0] = S90reg;
assign S91[LFSR_S-1:0] = S91reg;
assign S92[LFSR_S-1:0] = S92reg;
assign S93[LFSR_S-1:0] = S93reg;
assign S94[LFSR_S-1:0] = S94reg;
assign S95[LFSR_S-1:0] = S95reg;
assign S96[LFSR_S-1:0] = S96reg;
assign S97[LFSR_S-1:0] = S97reg;
assign S98[LFSR_S-1:0] = S98reg;
assign S99[LFSR_S-1:0] = S99reg;
assign S100[LFSR_S-1:0] = S100reg;
assign S101[LFSR_S-1:0] = S101reg;
assign S102[LFSR_S-1:0] = S102reg;
assign S103[LFSR_S-1:0] = S103reg;
assign S104[LFSR_S-1:0] = S104reg;
assign S105[LFSR_S-1:0] = S105reg;
assign S106[LFSR_S-1:0] = S106reg;
assign S107[LFSR_S-1:0] = S107reg;
assign S108[LFSR_S-1:0] = S108reg;
assign S109[LFSR_S-1:0] = S109reg;
assign S110[LFSR_S-1:0] = S110reg;
assign S111[LFSR_S-1:0] = S111reg;
assign S112[LFSR_S-1:0] = S112reg;
assign S113[LFSR_S-1:0] = S113reg;
assign S114[LFSR_S-1:0] = S114reg;
assign S115[LFSR_S-1:0] = S115reg;
assign S116[LFSR_S-1:0] = S116reg;
assign S117[LFSR_S-1:0] = S117reg;
assign S118[LFSR_S-1:0] = S118reg;
assign S119[LFSR_S-1:0] = S119reg;
assign S120[LFSR_S-1:0] = S120reg;
assign S121[LFSR_S-1:0] = S121reg;
assign S122[LFSR_S-1:0] = S122reg;
assign S123[LFSR_S-1:0] = S123reg;
assign S124[LFSR_S-1:0] = S124reg;
assign S125[LFSR_S-1:0] = S125reg;
assign S126[LFSR_S-1:0] = S126reg;
assign S127[LFSR_S-1:0] = S127reg;
assign S128[LFSR_S-1:0] = S128reg;
assign S129[LFSR_S-1:0] = S129reg;
assign S130[LFSR_S-1:0] = S130reg;
assign S131[LFSR_S-1:0] = S131reg;
assign S132[LFSR_S-1:0] = S132reg;
assign S133[LFSR_S-1:0] = S133reg;
assign S134[LFSR_S-1:0] = S134reg;
assign S135[LFSR_S-1:0] = S135reg;
assign S136[LFSR_S-1:0] = S136reg;
assign S137[LFSR_S-1:0] = S137reg;
assign S138[LFSR_S-1:0] = S138reg;
assign S139[LFSR_S-1:0] = S139reg;
assign S140[LFSR_S-1:0] = S140reg;
assign S141[LFSR_S-1:0] = S141reg;
assign S142[LFSR_S-1:0] = S142reg;
assign S143[LFSR_S-1:0] = S143reg;
assign S144[LFSR_S-1:0] = S144reg;
assign S145[LFSR_S-1:0] = S145reg;
assign S146[LFSR_S-1:0] = S146reg;
assign S147[LFSR_S-1:0] = S147reg;
assign S148[LFSR_S-1:0] = S148reg;
assign S149[LFSR_S-1:0] = S149reg;
assign S150[LFSR_S-1:0] = S150reg;
assign S151[LFSR_S-1:0] = S151reg;
assign S152[LFSR_S-1:0] = S152reg;
assign S153[LFSR_S-1:0] = S153reg;
assign S154[LFSR_S-1:0] = S154reg;
assign S155[LFSR_S-1:0] = S155reg;
assign S156[LFSR_S-1:0] = S156reg;
assign S157[LFSR_S-1:0] = S157reg;
assign S158[LFSR_S-1:0] = S158reg;
assign S159[LFSR_S-1:0] = S159reg;
assign S160[LFSR_S-1:0] = S160reg;
assign S161[LFSR_S-1:0] = S161reg;
assign S162[LFSR_S-1:0] = S162reg;
assign S163[LFSR_S-1:0] = S163reg;
assign S164[LFSR_S-1:0] = S164reg;
assign S165[LFSR_S-1:0] = S165reg;
assign S166[LFSR_S-1:0] = S166reg;
assign S167[LFSR_S-1:0] = S167reg;
assign S168[LFSR_S-1:0] = S168reg;
assign S169[LFSR_S-1:0] = S169reg;
assign S170[LFSR_S-1:0] = S170reg;
assign S171[LFSR_S-1:0] = S171reg;
assign S172[LFSR_S-1:0] = S172reg;
assign S173[LFSR_S-1:0] = S173reg;
assign S174[LFSR_S-1:0] = S174reg;
assign S175[LFSR_S-1:0] = S175reg;
assign S176[LFSR_S-1:0] = S176reg;
assign S177[LFSR_S-1:0] = S177reg;
assign S178[LFSR_S-1:0] = S178reg;
assign S179[LFSR_S-1:0] = S179reg;
assign S180[LFSR_S-1:0] = S180reg;
assign S181[LFSR_S-1:0] = S181reg;
assign S182[LFSR_S-1:0] = S182reg;
assign S183[LFSR_S-1:0] = S183reg;
assign S184[LFSR_S-1:0] = S184reg;
assign S185[LFSR_S-1:0] = S185reg;
assign S186[LFSR_S-1:0] = S186reg;
assign S187[LFSR_S-1:0] = S187reg;
assign S188[LFSR_S-1:0] = S188reg;
assign S189[LFSR_S-1:0] = S189reg;
assign S190[LFSR_S-1:0] = S190reg;
assign S191[LFSR_S-1:0] = S191reg;
assign S192[LFSR_S-1:0] = S192reg;
assign S193[LFSR_S-1:0] = S193reg;
assign S194[LFSR_S-1:0] = S194reg;
assign S195[LFSR_S-1:0] = S195reg;
assign S196[LFSR_S-1:0] = S196reg;
assign S197[LFSR_S-1:0] = S197reg;
assign S198[LFSR_S-1:0] = S198reg;
assign S199[LFSR_S-1:0] = S199reg;
assign S200[LFSR_S-1:0] = S200reg;
assign S201[LFSR_S-1:0] = S201reg;
assign S202[LFSR_S-1:0] = S202reg;
assign S203[LFSR_S-1:0] = S203reg;
assign S204[LFSR_S-1:0] = S204reg;
assign S205[LFSR_S-1:0] = S205reg;
assign S206[LFSR_S-1:0] = S206reg;
assign S207[LFSR_S-1:0] = S207reg;
assign S208[LFSR_S-1:0] = S208reg;
assign S209[LFSR_S-1:0] = S209reg;
assign S210[LFSR_S-1:0] = S210reg;
assign S211[LFSR_S-1:0] = S211reg;
assign S212[LFSR_S-1:0] = S212reg;
assign S213[LFSR_S-1:0] = S213reg;
assign S214[LFSR_S-1:0] = S214reg;
assign S215[LFSR_S-1:0] = S215reg;
assign S216[LFSR_S-1:0] = S216reg;
assign S217[LFSR_S-1:0] = S217reg;
assign S218[LFSR_S-1:0] = S218reg;
assign S219[LFSR_S-1:0] = S219reg;
assign S220[LFSR_S-1:0] = S220reg;
assign S221[LFSR_S-1:0] = S221reg;
assign S222[LFSR_S-1:0] = S222reg;
assign S223[LFSR_S-1:0] = S223reg;
assign S224[LFSR_S-1:0] = S224reg;
assign S225[LFSR_S-1:0] = S225reg;
assign S226[LFSR_S-1:0] = S226reg;
assign S227[LFSR_S-1:0] = S227reg;
assign S228[LFSR_S-1:0] = S228reg;
assign S229[LFSR_S-1:0] = S229reg;
assign S230[LFSR_S-1:0] = S230reg;
assign S231[LFSR_S-1:0] = S231reg;
assign S232[LFSR_S-1:0] = S232reg;
assign S233[LFSR_S-1:0] = S233reg;
assign S234[LFSR_S-1:0] = S234reg;
assign S235[LFSR_S-1:0] = S235reg;
assign S236[LFSR_S-1:0] = S236reg;
assign S237[LFSR_S-1:0] = S237reg;
assign S238[LFSR_S-1:0] = S238reg;
assign S239[LFSR_S-1:0] = S239reg;
assign S240[LFSR_S-1:0] = S240reg;
assign S241[LFSR_S-1:0] = S241reg;
assign S242[LFSR_S-1:0] = S242reg;
assign S243[LFSR_S-1:0] = S243reg;
assign S244[LFSR_S-1:0] = S244reg;
assign S245[LFSR_S-1:0] = S245reg;
assign S246[LFSR_S-1:0] = S246reg;
assign S247[LFSR_S-1:0] = S247reg;
assign S248[LFSR_S-1:0] = S248reg;
assign S249[LFSR_S-1:0] = S249reg;
assign S250[LFSR_S-1:0] = S250reg;
assign S251[LFSR_S-1:0] = S251reg;
assign S252[LFSR_S-1:0] = S252reg;
assign S253[LFSR_S-1:0] = S253reg;
assign S254[LFSR_S-1:0] = S254reg;
assign S255[LFSR_S-1:0] = S255reg;
assign S256[LFSR_S-1:0] = S256reg;
assign S257[LFSR_S-1:0] = S257reg;
assign S258[LFSR_S-1:0] = S258reg;
assign S259[LFSR_S-1:0] = S259reg;
assign S260[LFSR_S-1:0] = S260reg;
assign S261[LFSR_S-1:0] = S261reg;
assign S262[LFSR_S-1:0] = S262reg;
assign S263[LFSR_S-1:0] = S263reg;
assign S264[LFSR_S-1:0] = S264reg;
assign S265[LFSR_S-1:0] = S265reg;
assign S266[LFSR_S-1:0] = S266reg;
assign S267[LFSR_S-1:0] = S267reg;
assign S268[LFSR_S-1:0] = S268reg;
assign S269[LFSR_S-1:0] = S269reg;
assign S270[LFSR_S-1:0] = S270reg;
assign S271[LFSR_S-1:0] = S271reg;
assign S272[LFSR_S-1:0] = S272reg;
assign S273[LFSR_S-1:0] = S273reg;
assign S274[LFSR_S-1:0] = S274reg;
assign S275[LFSR_S-1:0] = S275reg;
assign S276[LFSR_S-1:0] = S276reg;
assign S277[LFSR_S-1:0] = S277reg;
assign S278[LFSR_S-1:0] = S278reg;
assign S279[LFSR_S-1:0] = S279reg;

always @(posedge INIT) begin

	if ((n1==4)&(ndiff!=4)) begin
		n1 = 1'b1;
		ndiff = ndiff + 1'b1;
	end
	else if (n1==4) begin
		n1 = 1'b1;
		ndiff = 1'b1;
	end
	else n1 = n1+1'b1;

	if (n1==1) n2 = ndiff;
	else if (n2==4) n2 = 1;
	else n2 = n2 + 1'b1;

	if (n1==1) begin
		S0reg [LFSR_S-1:0] <= 16'b1000000110001111;
		S1reg [LFSR_S-1:0] <= 16'b1001001010111111;
		S2reg [LFSR_S-1:0] <= 16'b0011001011010100;
		S3reg [LFSR_S-1:0] <= 16'b0110101011000110;
		S4reg [LFSR_S-1:0] <= 16'b0010110100110000;
		S5reg [LFSR_S-1:0] <= 16'b1110100110010000;
		S6reg [LFSR_S-1:0] <= 16'b1001110100011010;
		S7reg [LFSR_S-1:0] <= 16'b1001001111110111;
		S8reg [LFSR_S-1:0] <= 16'b1000111001101110;
		S9reg [LFSR_S-1:0] <= 16'b1110011111101011;
		S10reg [LFSR_S-1:0] <= 16'b0011100100001100;
		S11reg [LFSR_S-1:0] <= 16'b1001111100001111;
		S12reg [LFSR_S-1:0] <= 16'b0011111000111101;
		S13reg [LFSR_S-1:0] <= 16'b1110110110001101;
		S14reg [LFSR_S-1:0] <= 16'b1011010010110011;
		S15reg [LFSR_S-1:0] <= 16'b1010100000110010;
		S16reg [LFSR_S-1:0] <= 16'b0001000000111000;
		S17reg [LFSR_S-1:0] <= 16'b0100010101101100;
		S18reg [LFSR_S-1:0] <= 16'b1101110011110101;
		S19reg [LFSR_S-1:0] <= 16'b0100111010011000;
		S20reg [LFSR_S-1:0] <= 16'b1010101010101101;
		S21reg [LFSR_S-1:0] <= 16'b0101110011001110;
		S22reg [LFSR_S-1:0] <= 16'b0100101100001000;
		S23reg [LFSR_S-1:0] <= 16'b1010000100101010;
		S24reg [LFSR_S-1:0] <= 16'b1111101110010010;
		S25reg [LFSR_S-1:0] <= 16'b1110000010000000;
		S26reg [LFSR_S-1:0] <= 16'b1001101011011110;
		S27reg [LFSR_S-1:0] <= 16'b0001001100110111;
		S28reg [LFSR_S-1:0] <= 16'b1111011111100001;
		S29reg [LFSR_S-1:0] <= 16'b1011110011111001;
		S30reg [LFSR_S-1:0] <= 16'b1110010101011111;
		S31reg [LFSR_S-1:0] <= 16'b0011001100010111;
		S32reg [LFSR_S-1:0] <= 16'b0001010000010111;
		S33reg [LFSR_S-1:0] <= 16'b0100000110110011;
		S34reg [LFSR_S-1:0] <= 16'b1110100001001001;
		S35reg [LFSR_S-1:0] <= 16'b1101111000010000;
		S36reg [LFSR_S-1:0] <= 16'b0000010111111000;
		S37reg [LFSR_S-1:0] <= 16'b0101111111010011;
		S38reg [LFSR_S-1:0] <= 16'b1101001010010110;
		S39reg [LFSR_S-1:0] <= 16'b0001000110001000;
		S40reg [LFSR_S-1:0] <= 16'b0100000001101000;
		S41reg [LFSR_S-1:0] <= 16'b1110111111000101;
		S42reg [LFSR_S-1:0] <= 16'b1111000011111101;
		S43reg [LFSR_S-1:0] <= 16'b0111110111011110;
		S44reg [LFSR_S-1:0] <= 16'b0010110000100010;
		S45reg [LFSR_S-1:0] <= 16'b0101110111000010;
		S46reg [LFSR_S-1:0] <= 16'b1111110100011011;
		S47reg [LFSR_S-1:0] <= 16'b0101001100011101;
		S48reg [LFSR_S-1:0] <= 16'b1001110111111011;
		S49reg [LFSR_S-1:0] <= 16'b0000010000010010;
		S50reg [LFSR_S-1:0] <= 16'b1101011001111001;
		S51reg [LFSR_S-1:0] <= 16'b1011001101100111;
		S52reg [LFSR_S-1:0] <= 16'b1011100010001001;
		S53reg [LFSR_S-1:0] <= 16'b1111000010001111;
		S54reg [LFSR_S-1:0] <= 16'b0100011010101100;
		S55reg [LFSR_S-1:0] <= 16'b1000101110000101;
		S56reg [LFSR_S-1:0] <= 16'b1100100111100101;
		S57reg [LFSR_S-1:0] <= 16'b0001000001010000;
		S58reg [LFSR_S-1:0] <= 16'b0011011110011010;
		S59reg [LFSR_S-1:0] <= 16'b1001000011110001;
		S60reg [LFSR_S-1:0] <= 16'b0100001101101000;
		S61reg [LFSR_S-1:0] <= 16'b0000111010000011;
		S62reg [LFSR_S-1:0] <= 16'b1010101000001011;
		S63reg [LFSR_S-1:0] <= 16'b1111011110101011;
		S64reg [LFSR_S-1:0] <= 16'b1100000000000010;
		S65reg [LFSR_S-1:0] <= 16'b1000010010101001;
		S66reg [LFSR_S-1:0] <= 16'b0000101000011000;
		S67reg [LFSR_S-1:0] <= 16'b0110010010011010;
		S68reg [LFSR_S-1:0] <= 16'b1001101011101111;
		S69reg [LFSR_S-1:0] <= 16'b0100011001000110;
		S70reg [LFSR_S-1:0] <= 16'b0011111101111100;
		S71reg [LFSR_S-1:0] <= 16'b0111101110000101;
		S72reg [LFSR_S-1:0] <= 16'b0101000100001101;
		S73reg [LFSR_S-1:0] <= 16'b0110100101111011;
		S74reg [LFSR_S-1:0] <= 16'b1011110110011011;
		S75reg [LFSR_S-1:0] <= 16'b0110010101111010;
		S76reg [LFSR_S-1:0] <= 16'b0000001101101000;
		S77reg [LFSR_S-1:0] <= 16'b1111100111011000;
		S78reg [LFSR_S-1:0] <= 16'b1010110001000010;
		S79reg [LFSR_S-1:0] <= 16'b0100110000110100;
		S80reg [LFSR_S-1:0] <= 16'b0010011011010001;
		S81reg [LFSR_S-1:0] <= 16'b1001000000101100;
		S82reg [LFSR_S-1:0] <= 16'b1010101100111101;
		S83reg [LFSR_S-1:0] <= 16'b1001010011011111;
		S84reg [LFSR_S-1:0] <= 16'b1010101110000000;
		S85reg [LFSR_S-1:0] <= 16'b1011110010010101;
		S86reg [LFSR_S-1:0] <= 16'b0101101111111100;
		S87reg [LFSR_S-1:0] <= 16'b1110010111110000;
		S88reg [LFSR_S-1:0] <= 16'b0101111101100110;
		S89reg [LFSR_S-1:0] <= 16'b0101101010001011;
		S90reg [LFSR_S-1:0] <= 16'b1100001001001101;
		S91reg [LFSR_S-1:0] <= 16'b0000101011010011;
		S92reg [LFSR_S-1:0] <= 16'b1000100000011100;
		S93reg [LFSR_S-1:0] <= 16'b1011010101001010;
		S94reg [LFSR_S-1:0] <= 16'b1110100100110101;
		S95reg [LFSR_S-1:0] <= 16'b0100111110000010;
		S96reg [LFSR_S-1:0] <= 16'b1000001100100101;
		S97reg [LFSR_S-1:0] <= 16'b1011011001100000;
		S98reg [LFSR_S-1:0] <= 16'b0011101010101101;
		S99reg [LFSR_S-1:0] <= 16'b0000000000001010;
		S100reg [LFSR_S-1:0] <= 16'b0100011010011111;
		S101reg [LFSR_S-1:0] <= 16'b0111010101101101;
		S102reg [LFSR_S-1:0] <= 16'b0111101010101000;
		S103reg [LFSR_S-1:0] <= 16'b0100010101100000;
		S104reg [LFSR_S-1:0] <= 16'b1110110001011111;
		S105reg [LFSR_S-1:0] <= 16'b0001111100111111;
		S106reg [LFSR_S-1:0] <= 16'b0111000101001011;
		S107reg [LFSR_S-1:0] <= 16'b1111000111101011;
		S108reg [LFSR_S-1:0] <= 16'b1011010011100101;
		S109reg [LFSR_S-1:0] <= 16'b1011111111100011;
		S110reg [LFSR_S-1:0] <= 16'b1011011110011111;
		S111reg [LFSR_S-1:0] <= 16'b0101100001010101;
		S112reg [LFSR_S-1:0] <= 16'b0101011010011011;
		S113reg [LFSR_S-1:0] <= 16'b1111100110110101;
		S114reg [LFSR_S-1:0] <= 16'b0101111000001001;
		S115reg [LFSR_S-1:0] <= 16'b1011100010011001;
		S116reg [LFSR_S-1:0] <= 16'b1111010001100110;
		S117reg [LFSR_S-1:0] <= 16'b1111110010111111;
		S118reg [LFSR_S-1:0] <= 16'b1000001101111011;
		S119reg [LFSR_S-1:0] <= 16'b0110010110000111;
		S120reg [LFSR_S-1:0] <= 16'b0001110110010001;
		S121reg [LFSR_S-1:0] <= 16'b0110100010101000;
		S122reg [LFSR_S-1:0] <= 16'b0001110001010110;
		S123reg [LFSR_S-1:0] <= 16'b0010001011010100;
		S124reg [LFSR_S-1:0] <= 16'b1101011011101101;
		S125reg [LFSR_S-1:0] <= 16'b0111101001010000;
		S126reg [LFSR_S-1:0] <= 16'b0111001110100111;
		S127reg [LFSR_S-1:0] <= 16'b1001110111001000;
		S128reg [LFSR_S-1:0] <= 16'b0101001010001000;
		S129reg [LFSR_S-1:0] <= 16'b1010011001111001;
		S130reg [LFSR_S-1:0] <= 16'b0011000110110010;
		S131reg [LFSR_S-1:0] <= 16'b1010000001010101;
		S132reg [LFSR_S-1:0] <= 16'b1010100000000011;
		S133reg [LFSR_S-1:0] <= 16'b0101001111100110;
		S134reg [LFSR_S-1:0] <= 16'b0101111110001010;
		S135reg [LFSR_S-1:0] <= 16'b0100010100101000;
		S136reg [LFSR_S-1:0] <= 16'b0110101101010001;
		S137reg [LFSR_S-1:0] <= 16'b0001011010101110;
		S138reg [LFSR_S-1:0] <= 16'b1000001001100001;
		S139reg [LFSR_S-1:0] <= 16'b1100111011100011;
	end
	if (n2==1) begin
		S140reg [LFSR_S-1:0] <= 16'b1001100011110000;
		S141reg [LFSR_S-1:0] <= 16'b1100100011000111;
		S142reg [LFSR_S-1:0] <= 16'b0101101101010010;
		S143reg [LFSR_S-1:0] <= 16'b0000100000111000;
		S144reg [LFSR_S-1:0] <= 16'b0111001101111101;
		S145reg [LFSR_S-1:0] <= 16'b1000001010110111;
		S146reg [LFSR_S-1:0] <= 16'b1101100011011001;
		S147reg [LFSR_S-1:0] <= 16'b0000101111101010;
		S148reg [LFSR_S-1:0] <= 16'b1000111100111111;
		S149reg [LFSR_S-1:0] <= 16'b0011001000101000;
		S150reg [LFSR_S-1:0] <= 16'b0001011011110101;
		S151reg [LFSR_S-1:0] <= 16'b1100100010101011;
		S152reg [LFSR_S-1:0] <= 16'b1110110001110101;
		S153reg [LFSR_S-1:0] <= 16'b1010111110100100;
		S154reg [LFSR_S-1:0] <= 16'b0010011100111111;
		S155reg [LFSR_S-1:0] <= 16'b0001001110010111;
		S156reg [LFSR_S-1:0] <= 16'b0001100011010100;
		S157reg [LFSR_S-1:0] <= 16'b1000100001001101;
		S158reg [LFSR_S-1:0] <= 16'b1011010000100011;
		S159reg [LFSR_S-1:0] <= 16'b1001000111000001;
		S160reg [LFSR_S-1:0] <= 16'b0011010010100010;
		S161reg [LFSR_S-1:0] <= 16'b1000100101110011;
		S162reg [LFSR_S-1:0] <= 16'b1011001100000001;
		S163reg [LFSR_S-1:0] <= 16'b0101011001111101;
		S164reg [LFSR_S-1:0] <= 16'b0011011100000001;
		S165reg [LFSR_S-1:0] <= 16'b0101000101000100;
		S166reg [LFSR_S-1:0] <= 16'b0110111101001010;
		S167reg [LFSR_S-1:0] <= 16'b0010001000101000;
		S168reg [LFSR_S-1:0] <= 16'b0011010111100110;
		S169reg [LFSR_S-1:0] <= 16'b0111011111110011;
		S170reg [LFSR_S-1:0] <= 16'b0010001111011110;
		S171reg [LFSR_S-1:0] <= 16'b1111010111011101;
		S172reg [LFSR_S-1:0] <= 16'b1010110100011001;
		S173reg [LFSR_S-1:0] <= 16'b1011101100010001;
		S174reg [LFSR_S-1:0] <= 16'b0100001101110010;
		S175reg [LFSR_S-1:0] <= 16'b1001100000011110;
		S176reg [LFSR_S-1:0] <= 16'b0010111100110110;
		S177reg [LFSR_S-1:0] <= 16'b0100010101000100;
		S178reg [LFSR_S-1:0] <= 16'b1100101010001001;
		S179reg [LFSR_S-1:0] <= 16'b1111100101101101;
		S180reg [LFSR_S-1:0] <= 16'b0111110111001010;
		S181reg [LFSR_S-1:0] <= 16'b0010110010110110;
		S182reg [LFSR_S-1:0] <= 16'b0100100111100100;
		S183reg [LFSR_S-1:0] <= 16'b1101101000111011;
		S184reg [LFSR_S-1:0] <= 16'b1110011001110011;
		S185reg [LFSR_S-1:0] <= 16'b0101111100110000;
		S186reg [LFSR_S-1:0] <= 16'b1111100101100001;
		S187reg [LFSR_S-1:0] <= 16'b1100101010111100;
		S188reg [LFSR_S-1:0] <= 16'b1101101011001111;
		S189reg [LFSR_S-1:0] <= 16'b0101111111111101;
		S190reg [LFSR_S-1:0] <= 16'b1111011100111111;
		S191reg [LFSR_S-1:0] <= 16'b1100100011100100;
		S192reg [LFSR_S-1:0] <= 16'b0001110010011101;
		S193reg [LFSR_S-1:0] <= 16'b0110110100111010;
		S194reg [LFSR_S-1:0] <= 16'b1100000001111111;
		S195reg [LFSR_S-1:0] <= 16'b0111100001100010;
		S196reg [LFSR_S-1:0] <= 16'b0011010010110001;
		S197reg [LFSR_S-1:0] <= 16'b1111101111110001;
		S198reg [LFSR_S-1:0] <= 16'b1011100110111001;
		S199reg [LFSR_S-1:0] <= 16'b0100000000111000;
		S200reg [LFSR_S-1:0] <= 16'b0001011110110111;
		S201reg [LFSR_S-1:0] <= 16'b1000000100011010;
		S202reg [LFSR_S-1:0] <= 16'b1011000110101101;
		S203reg [LFSR_S-1:0] <= 16'b1011001010100011;
		S204reg [LFSR_S-1:0] <= 16'b0111101101011110;
		S205reg [LFSR_S-1:0] <= 16'b0110110101110101;
		S206reg [LFSR_S-1:0] <= 16'b0000110011000100;
		S207reg [LFSR_S-1:0] <= 16'b0111100001101101;
		S208reg [LFSR_S-1:0] <= 16'b0011001010110101;
		S209reg [LFSR_S-1:0] <= 16'b0010111010011100;
		S210reg [LFSR_S-1:0] <= 16'b0001010101110110;
		S211reg [LFSR_S-1:0] <= 16'b1110111001001011;
		S212reg [LFSR_S-1:0] <= 16'b1110111100110011;
		S213reg [LFSR_S-1:0] <= 16'b0110111111100100;
		S214reg [LFSR_S-1:0] <= 16'b1000001001100001;
		S215reg [LFSR_S-1:0] <= 16'b1001011100001001;
		S216reg [LFSR_S-1:0] <= 16'b0010001011101100;
		S217reg [LFSR_S-1:0] <= 16'b1010100110111001;
		S218reg [LFSR_S-1:0] <= 16'b0110011101110010;
		S219reg [LFSR_S-1:0] <= 16'b1010111001110111;
		S220reg [LFSR_S-1:0] <= 16'b0001001000000110;
		S221reg [LFSR_S-1:0] <= 16'b1011010100010001;
		S222reg [LFSR_S-1:0] <= 16'b0110100110101011;
		S223reg [LFSR_S-1:0] <= 16'b1110100001011100;
		S224reg [LFSR_S-1:0] <= 16'b1101010100000001;
		S225reg [LFSR_S-1:0] <= 16'b0011010101010100;
		S226reg [LFSR_S-1:0] <= 16'b0010001111010100;
		S227reg [LFSR_S-1:0] <= 16'b1001000000110111;
		S228reg [LFSR_S-1:0] <= 16'b0001000001001100;
		S229reg [LFSR_S-1:0] <= 16'b1010010110101011;
		S230reg [LFSR_S-1:0] <= 16'b0000010000010100;
		S231reg [LFSR_S-1:0] <= 16'b1111100100001011;
		S232reg [LFSR_S-1:0] <= 16'b1010110101000011;
		S233reg [LFSR_S-1:0] <= 16'b1110110010100010;
		S234reg [LFSR_S-1:0] <= 16'b0000111001100100;
		S235reg [LFSR_S-1:0] <= 16'b0010100001000000;
		S236reg [LFSR_S-1:0] <= 16'b1010101010100111;
		S237reg [LFSR_S-1:0] <= 16'b0010100100010100;
		S238reg [LFSR_S-1:0] <= 16'b0010101011100101;
		S239reg [LFSR_S-1:0] <= 16'b0110101111111110;
		S240reg [LFSR_S-1:0] <= 16'b0010101111011111;
		S241reg [LFSR_S-1:0] <= 16'b0010110101011000;
		S242reg [LFSR_S-1:0] <= 16'b0000001101110010;
		S243reg [LFSR_S-1:0] <= 16'b1100111010000001;
		S244reg [LFSR_S-1:0] <= 16'b1011001001001111;
		S245reg [LFSR_S-1:0] <= 16'b1000000110000110;
		S246reg [LFSR_S-1:0] <= 16'b1100110000101000;
		S247reg [LFSR_S-1:0] <= 16'b0001101100110100;
		S248reg [LFSR_S-1:0] <= 16'b0010111111001010;
		S249reg [LFSR_S-1:0] <= 16'b1111001000001001;
		S250reg [LFSR_S-1:0] <= 16'b1111101000001001;
		S251reg [LFSR_S-1:0] <= 16'b0010101100100001;
		S252reg [LFSR_S-1:0] <= 16'b1100000101000010;
		S253reg [LFSR_S-1:0] <= 16'b1000010001001101;
		S254reg [LFSR_S-1:0] <= 16'b0100000110001001;
		S255reg [LFSR_S-1:0] <= 16'b1001011000011010;
		S256reg [LFSR_S-1:0] <= 16'b0001000011010011;
		S257reg [LFSR_S-1:0] <= 16'b0001010111110100;
		S258reg [LFSR_S-1:0] <= 16'b0101000010101110;
		S259reg [LFSR_S-1:0] <= 16'b0111100000011111;
		S260reg [LFSR_S-1:0] <= 16'b1010000100101010;
		S261reg [LFSR_S-1:0] <= 16'b0101111110100001;
		S262reg [LFSR_S-1:0] <= 16'b1100010010101010;
		S263reg [LFSR_S-1:0] <= 16'b1000110011000010;
		S264reg [LFSR_S-1:0] <= 16'b0000011111111100;
		S265reg [LFSR_S-1:0] <= 16'b0101100101110111;
		S266reg [LFSR_S-1:0] <= 16'b0110100100010010;
		S267reg [LFSR_S-1:0] <= 16'b1100110101110100;
		S268reg [LFSR_S-1:0] <= 16'b1010010011100011;
		S269reg [LFSR_S-1:0] <= 16'b0101011011010000;
		S270reg [LFSR_S-1:0] <= 16'b0001011000101010;
		S271reg [LFSR_S-1:0] <= 16'b0000001101011000;
		S272reg [LFSR_S-1:0] <= 16'b1010000111101011;
		S273reg [LFSR_S-1:0] <= 16'b1101001011011010;
		S274reg [LFSR_S-1:0] <= 16'b0100101001000000;
		S275reg [LFSR_S-1:0] <= 16'b1100011100101101;
		S276reg [LFSR_S-1:0] <= 16'b1110100011001110;
		S277reg [LFSR_S-1:0] <= 16'b0101111000001100;
		S278reg [LFSR_S-1:0] <= 16'b0110011111111100;
		S279reg [LFSR_S-1:0] <= 16'b0010101001010100;
	end
	if (n1==2) begin
		S0reg [LFSR_S-1:0] <= 16'b1110001100000101;
		S1reg [LFSR_S-1:0] <= 16'b1111000000111100;
		S2reg [LFSR_S-1:0] <= 16'b0000001010110110;
		S3reg [LFSR_S-1:0] <= 16'b1000100000001111;
		S4reg [LFSR_S-1:0] <= 16'b1111010011010011;
		S5reg [LFSR_S-1:0] <= 16'b1010011010101001;
		S6reg [LFSR_S-1:0] <= 16'b1000110010011100;
		S7reg [LFSR_S-1:0] <= 16'b0111100101010111;
		S8reg [LFSR_S-1:0] <= 16'b0110001010000010;
		S9reg [LFSR_S-1:0] <= 16'b1010100010111100;
		S10reg [LFSR_S-1:0] <= 16'b0010001010001000;
		S11reg [LFSR_S-1:0] <= 16'b1110000001110111;
		S12reg [LFSR_S-1:0] <= 16'b1101100000011001;
		S13reg [LFSR_S-1:0] <= 16'b1010110100000011;
		S14reg [LFSR_S-1:0] <= 16'b1010011101111011;
		S15reg [LFSR_S-1:0] <= 16'b0101001010111100;
		S16reg [LFSR_S-1:0] <= 16'b1000110010101010;
		S17reg [LFSR_S-1:0] <= 16'b0100100001100010;
		S18reg [LFSR_S-1:0] <= 16'b1110110100101001;
		S19reg [LFSR_S-1:0] <= 16'b0010011011000011;
		S20reg [LFSR_S-1:0] <= 16'b1110011100100101;
		S21reg [LFSR_S-1:0] <= 16'b1011010100100101;
		S22reg [LFSR_S-1:0] <= 16'b0100101010001011;
		S23reg [LFSR_S-1:0] <= 16'b1111011101001001;
		S24reg [LFSR_S-1:0] <= 16'b1001100001110011;
		S25reg [LFSR_S-1:0] <= 16'b1111111111110111;
		S26reg [LFSR_S-1:0] <= 16'b0100101111000010;
		S27reg [LFSR_S-1:0] <= 16'b1010010000111101;
		S28reg [LFSR_S-1:0] <= 16'b0111010100100010;
		S29reg [LFSR_S-1:0] <= 16'b1001111000000110;
		S30reg [LFSR_S-1:0] <= 16'b1010010000100111;
		S31reg [LFSR_S-1:0] <= 16'b1111100110111111;
		S32reg [LFSR_S-1:0] <= 16'b0001000000011000;
		S33reg [LFSR_S-1:0] <= 16'b1000110010111101;
		S34reg [LFSR_S-1:0] <= 16'b1001010011111111;
		S35reg [LFSR_S-1:0] <= 16'b0100010110110000;
		S36reg [LFSR_S-1:0] <= 16'b1100111000111110;
		S37reg [LFSR_S-1:0] <= 16'b1111110011100001;
		S38reg [LFSR_S-1:0] <= 16'b1010110010001110;
		S39reg [LFSR_S-1:0] <= 16'b0011011011110001;
		S40reg [LFSR_S-1:0] <= 16'b1000111100101101;
		S41reg [LFSR_S-1:0] <= 16'b1101100110110011;
		S42reg [LFSR_S-1:0] <= 16'b0011011101011011;
		S43reg [LFSR_S-1:0] <= 16'b0010011001110100;
		S44reg [LFSR_S-1:0] <= 16'b1101110010100001;
		S45reg [LFSR_S-1:0] <= 16'b1101110111101101;
		S46reg [LFSR_S-1:0] <= 16'b0110101110000110;
		S47reg [LFSR_S-1:0] <= 16'b1111111010100010;
		S48reg [LFSR_S-1:0] <= 16'b0010111000000100;
		S49reg [LFSR_S-1:0] <= 16'b1111010000100000;
		S50reg [LFSR_S-1:0] <= 16'b0011010100010101;
		S51reg [LFSR_S-1:0] <= 16'b1010010001010111;
		S52reg [LFSR_S-1:0] <= 16'b1110100110110011;
		S53reg [LFSR_S-1:0] <= 16'b0001110001000000;
		S54reg [LFSR_S-1:0] <= 16'b0001000001011000;
		S55reg [LFSR_S-1:0] <= 16'b1001111101011110;
		S56reg [LFSR_S-1:0] <= 16'b1111100011100101;
		S57reg [LFSR_S-1:0] <= 16'b0001001111101101;
		S58reg [LFSR_S-1:0] <= 16'b1101110010010011;
		S59reg [LFSR_S-1:0] <= 16'b0010000000110110;
		S60reg [LFSR_S-1:0] <= 16'b0110110010100001;
		S61reg [LFSR_S-1:0] <= 16'b1001100110010100;
		S62reg [LFSR_S-1:0] <= 16'b0000111000111000;
		S63reg [LFSR_S-1:0] <= 16'b0000011011010010;
		S64reg [LFSR_S-1:0] <= 16'b0110001011011000;
		S65reg [LFSR_S-1:0] <= 16'b1111110010110101;
		S66reg [LFSR_S-1:0] <= 16'b1100011110010101;
		S67reg [LFSR_S-1:0] <= 16'b1011010001110100;
		S68reg [LFSR_S-1:0] <= 16'b1101100011110011;
		S69reg [LFSR_S-1:0] <= 16'b1100100111110111;
		S70reg [LFSR_S-1:0] <= 16'b1010111111011001;
		S71reg [LFSR_S-1:0] <= 16'b0111010001110100;
		S72reg [LFSR_S-1:0] <= 16'b1111001011111011;
		S73reg [LFSR_S-1:0] <= 16'b1000101011110100;
		S74reg [LFSR_S-1:0] <= 16'b1011001100011100;
		S75reg [LFSR_S-1:0] <= 16'b1110010000110100;
		S76reg [LFSR_S-1:0] <= 16'b0011001100111010;
		S77reg [LFSR_S-1:0] <= 16'b0001101100111100;
		S78reg [LFSR_S-1:0] <= 16'b1010110110100011;
		S79reg [LFSR_S-1:0] <= 16'b1110011111001101;
		S80reg [LFSR_S-1:0] <= 16'b0100010110010010;
		S81reg [LFSR_S-1:0] <= 16'b0010101100100000;
		S82reg [LFSR_S-1:0] <= 16'b1010010010110110;
		S83reg [LFSR_S-1:0] <= 16'b1111001111100011;
		S84reg [LFSR_S-1:0] <= 16'b1111100001111100;
		S85reg [LFSR_S-1:0] <= 16'b0111011110010110;
		S86reg [LFSR_S-1:0] <= 16'b0001000011111000;
		S87reg [LFSR_S-1:0] <= 16'b0010000101110001;
		S88reg [LFSR_S-1:0] <= 16'b0000101110011001;
		S89reg [LFSR_S-1:0] <= 16'b1001100101110101;
		S90reg [LFSR_S-1:0] <= 16'b1000010000111010;
		S91reg [LFSR_S-1:0] <= 16'b0111110001011110;
		S92reg [LFSR_S-1:0] <= 16'b1100010101100100;
		S93reg [LFSR_S-1:0] <= 16'b0110011111000101;
		S94reg [LFSR_S-1:0] <= 16'b1001011001110011;
		S95reg [LFSR_S-1:0] <= 16'b0001010110000100;
		S96reg [LFSR_S-1:0] <= 16'b1001010001111010;
		S97reg [LFSR_S-1:0] <= 16'b1000101111001011;
		S98reg [LFSR_S-1:0] <= 16'b0110000111100111;
		S99reg [LFSR_S-1:0] <= 16'b0101001010010101;
		S100reg [LFSR_S-1:0] <= 16'b0011011000001111;
		S101reg [LFSR_S-1:0] <= 16'b1011110110001011;
		S102reg [LFSR_S-1:0] <= 16'b0001011110011000;
		S103reg [LFSR_S-1:0] <= 16'b1001011011011011;
		S104reg [LFSR_S-1:0] <= 16'b1010110010000110;
		S105reg [LFSR_S-1:0] <= 16'b0010000011100110;
		S106reg [LFSR_S-1:0] <= 16'b1001011101110111;
		S107reg [LFSR_S-1:0] <= 16'b1001100000001111;
		S108reg [LFSR_S-1:0] <= 16'b1010111100000101;
		S109reg [LFSR_S-1:0] <= 16'b1001111011111000;
		S110reg [LFSR_S-1:0] <= 16'b0000011011101010;
		S111reg [LFSR_S-1:0] <= 16'b1000101110111101;
		S112reg [LFSR_S-1:0] <= 16'b0001100100110110;
		S113reg [LFSR_S-1:0] <= 16'b1000101010110000;
		S114reg [LFSR_S-1:0] <= 16'b1011000010110011;
		S115reg [LFSR_S-1:0] <= 16'b0001010111111101;
		S116reg [LFSR_S-1:0] <= 16'b1000110101110010;
		S117reg [LFSR_S-1:0] <= 16'b1001010110000000;
		S118reg [LFSR_S-1:0] <= 16'b0100101001001101;
		S119reg [LFSR_S-1:0] <= 16'b1000110011101101;
		S120reg [LFSR_S-1:0] <= 16'b0110100011110111;
		S121reg [LFSR_S-1:0] <= 16'b1011101111000011;
		S122reg [LFSR_S-1:0] <= 16'b0000100100001000;
		S123reg [LFSR_S-1:0] <= 16'b0000001000110000;
		S124reg [LFSR_S-1:0] <= 16'b0101010000000000;
		S125reg [LFSR_S-1:0] <= 16'b0000001001100110;
		S126reg [LFSR_S-1:0] <= 16'b1010100101010010;
		S127reg [LFSR_S-1:0] <= 16'b1110001111110111;
		S128reg [LFSR_S-1:0] <= 16'b0011011000110100;
		S129reg [LFSR_S-1:0] <= 16'b1000010011101111;
		S130reg [LFSR_S-1:0] <= 16'b1101000000010101;
		S131reg [LFSR_S-1:0] <= 16'b1110111110111111;
		S132reg [LFSR_S-1:0] <= 16'b1111101101001001;
		S133reg [LFSR_S-1:0] <= 16'b0101010010001010;
		S134reg [LFSR_S-1:0] <= 16'b1010011101110000;
		S135reg [LFSR_S-1:0] <= 16'b0100111110111000;
		S136reg [LFSR_S-1:0] <= 16'b0000000001001100;
		S137reg [LFSR_S-1:0] <= 16'b1101010100111010;
		S138reg [LFSR_S-1:0] <= 16'b0100110111100110;
		S139reg [LFSR_S-1:0] <= 16'b0001110001101100;
	end
	if (n2==2) begin
		S140reg [LFSR_S-1:0] <= 16'b1010011001000100;
		S141reg [LFSR_S-1:0] <= 16'b1110010101010110;
		S142reg [LFSR_S-1:0] <= 16'b0101111001100010;
		S143reg [LFSR_S-1:0] <= 16'b0100000110110100;
		S144reg [LFSR_S-1:0] <= 16'b0111010110100010;
		S145reg [LFSR_S-1:0] <= 16'b1111111000110011;
		S146reg [LFSR_S-1:0] <= 16'b0111010111010010;
		S147reg [LFSR_S-1:0] <= 16'b0100010001000010;
		S148reg [LFSR_S-1:0] <= 16'b0010100111010011;
		S149reg [LFSR_S-1:0] <= 16'b0111110001100100;
		S150reg [LFSR_S-1:0] <= 16'b1100110100000101;
		S151reg [LFSR_S-1:0] <= 16'b1111110100100001;
		S152reg [LFSR_S-1:0] <= 16'b1001100011111011;
		S153reg [LFSR_S-1:0] <= 16'b0111011011010010;
		S154reg [LFSR_S-1:0] <= 16'b0010101001011010;
		S155reg [LFSR_S-1:0] <= 16'b0000101100100100;
		S156reg [LFSR_S-1:0] <= 16'b1001100111101101;
		S157reg [LFSR_S-1:0] <= 16'b1011010100111101;
		S158reg [LFSR_S-1:0] <= 16'b0000100011000010;
		S159reg [LFSR_S-1:0] <= 16'b1001111110100000;
		S160reg [LFSR_S-1:0] <= 16'b0100111101010111;
		S161reg [LFSR_S-1:0] <= 16'b1001010110001111;
		S162reg [LFSR_S-1:0] <= 16'b1010111001001010;
		S163reg [LFSR_S-1:0] <= 16'b0001100110100100;
		S164reg [LFSR_S-1:0] <= 16'b1010111100101110;
		S165reg [LFSR_S-1:0] <= 16'b0001100001110100;
		S166reg [LFSR_S-1:0] <= 16'b0101111111000111;
		S167reg [LFSR_S-1:0] <= 16'b1000101100110100;
		S168reg [LFSR_S-1:0] <= 16'b1011111111110101;
		S169reg [LFSR_S-1:0] <= 16'b1000100111011101;
		S170reg [LFSR_S-1:0] <= 16'b1001100001111011;
		S171reg [LFSR_S-1:0] <= 16'b0101110000000100;
		S172reg [LFSR_S-1:0] <= 16'b1011010010110101;
		S173reg [LFSR_S-1:0] <= 16'b0100111001000100;
		S174reg [LFSR_S-1:0] <= 16'b0111100110100101;
		S175reg [LFSR_S-1:0] <= 16'b1000111010111010;
		S176reg [LFSR_S-1:0] <= 16'b1101101110101001;
		S177reg [LFSR_S-1:0] <= 16'b1100010001101110;
		S178reg [LFSR_S-1:0] <= 16'b1001000100011001;
		S179reg [LFSR_S-1:0] <= 16'b0010101111010000;
		S180reg [LFSR_S-1:0] <= 16'b0100010011011011;
		S181reg [LFSR_S-1:0] <= 16'b0110000010101100;
		S182reg [LFSR_S-1:0] <= 16'b1110001111111101;
		S183reg [LFSR_S-1:0] <= 16'b1101010010011111;
		S184reg [LFSR_S-1:0] <= 16'b1100010111111000;
		S185reg [LFSR_S-1:0] <= 16'b0011010001101110;
		S186reg [LFSR_S-1:0] <= 16'b1110111100000010;
		S187reg [LFSR_S-1:0] <= 16'b0010010010000100;
		S188reg [LFSR_S-1:0] <= 16'b0100110111100110;
		S189reg [LFSR_S-1:0] <= 16'b1001101111110110;
		S190reg [LFSR_S-1:0] <= 16'b0110001111010101;
		S191reg [LFSR_S-1:0] <= 16'b0101000100100010;
		S192reg [LFSR_S-1:0] <= 16'b0000001000000010;
		S193reg [LFSR_S-1:0] <= 16'b1100011011111001;
		S194reg [LFSR_S-1:0] <= 16'b0111011101010101;
		S195reg [LFSR_S-1:0] <= 16'b0111101110010010;
		S196reg [LFSR_S-1:0] <= 16'b0011001101111101;
		S197reg [LFSR_S-1:0] <= 16'b0011101110110101;
		S198reg [LFSR_S-1:0] <= 16'b0010001010100000;
		S199reg [LFSR_S-1:0] <= 16'b0111100011101111;
		S200reg [LFSR_S-1:0] <= 16'b0010001001111010;
		S201reg [LFSR_S-1:0] <= 16'b1000100100010011;
		S202reg [LFSR_S-1:0] <= 16'b1011010111110110;
		S203reg [LFSR_S-1:0] <= 16'b0011110010101110;
		S204reg [LFSR_S-1:0] <= 16'b1100110001111110;
		S205reg [LFSR_S-1:0] <= 16'b0010110100001000;
		S206reg [LFSR_S-1:0] <= 16'b1000011011010011;
		S207reg [LFSR_S-1:0] <= 16'b0111000111010110;
		S208reg [LFSR_S-1:0] <= 16'b1101011100100111;
		S209reg [LFSR_S-1:0] <= 16'b0010011001100000;
		S210reg [LFSR_S-1:0] <= 16'b0101011001010111;
		S211reg [LFSR_S-1:0] <= 16'b1010110100110101;
		S212reg [LFSR_S-1:0] <= 16'b1000111011001000;
		S213reg [LFSR_S-1:0] <= 16'b1111010001100110;
		S214reg [LFSR_S-1:0] <= 16'b1001000101001101;
		S215reg [LFSR_S-1:0] <= 16'b0100101100110111;
		S216reg [LFSR_S-1:0] <= 16'b1111001010001011;
		S217reg [LFSR_S-1:0] <= 16'b0101001000101010;
		S218reg [LFSR_S-1:0] <= 16'b0001110110000010;
		S219reg [LFSR_S-1:0] <= 16'b0010101010000110;
		S220reg [LFSR_S-1:0] <= 16'b0000010101110110;
		S221reg [LFSR_S-1:0] <= 16'b1000000010101000;
		S222reg [LFSR_S-1:0] <= 16'b1100110010110011;
		S223reg [LFSR_S-1:0] <= 16'b1000101110000011;
		S224reg [LFSR_S-1:0] <= 16'b0110000010111100;
		S225reg [LFSR_S-1:0] <= 16'b1101111111010000;
		S226reg [LFSR_S-1:0] <= 16'b1100101111000011;
		S227reg [LFSR_S-1:0] <= 16'b0011010011000010;
		S228reg [LFSR_S-1:0] <= 16'b0000000011101100;
		S229reg [LFSR_S-1:0] <= 16'b0011000010000000;
		S230reg [LFSR_S-1:0] <= 16'b1110111110010011;
		S231reg [LFSR_S-1:0] <= 16'b0001001010101110;
		S232reg [LFSR_S-1:0] <= 16'b0010010110001010;
		S233reg [LFSR_S-1:0] <= 16'b0011011100110010;
		S234reg [LFSR_S-1:0] <= 16'b0001111010001010;
		S235reg [LFSR_S-1:0] <= 16'b0100111111111001;
		S236reg [LFSR_S-1:0] <= 16'b0000111100000110;
		S237reg [LFSR_S-1:0] <= 16'b0010000000101000;
		S238reg [LFSR_S-1:0] <= 16'b1011001100001111;
		S239reg [LFSR_S-1:0] <= 16'b1010111001010001;
		S240reg [LFSR_S-1:0] <= 16'b0001100110100010;
		S241reg [LFSR_S-1:0] <= 16'b1101110111110000;
		S242reg [LFSR_S-1:0] <= 16'b1100111100011001;
		S243reg [LFSR_S-1:0] <= 16'b0001101100010001;
		S244reg [LFSR_S-1:0] <= 16'b1101110100101110;
		S245reg [LFSR_S-1:0] <= 16'b1110010001100011;
		S246reg [LFSR_S-1:0] <= 16'b0100111000101110;
		S247reg [LFSR_S-1:0] <= 16'b1000011110001011;
		S248reg [LFSR_S-1:0] <= 16'b0000010110010111;
		S249reg [LFSR_S-1:0] <= 16'b0101101001010010;
		S250reg [LFSR_S-1:0] <= 16'b1001101110011111;
		S251reg [LFSR_S-1:0] <= 16'b0100110000110111;
		S252reg [LFSR_S-1:0] <= 16'b0001001000011100;
		S253reg [LFSR_S-1:0] <= 16'b0010011111011011;
		S254reg [LFSR_S-1:0] <= 16'b0101110111001001;
		S255reg [LFSR_S-1:0] <= 16'b1011001011101011;
		S256reg [LFSR_S-1:0] <= 16'b1010110010111101;
		S257reg [LFSR_S-1:0] <= 16'b0010111111100110;
		S258reg [LFSR_S-1:0] <= 16'b0110111001101010;
		S259reg [LFSR_S-1:0] <= 16'b1011001010101101;
		S260reg [LFSR_S-1:0] <= 16'b1101111100010011;
		S261reg [LFSR_S-1:0] <= 16'b1100100100100100;
		S262reg [LFSR_S-1:0] <= 16'b1110001100100011;
		S263reg [LFSR_S-1:0] <= 16'b1101110110011001;
		S264reg [LFSR_S-1:0] <= 16'b0101000000000100;
		S265reg [LFSR_S-1:0] <= 16'b0111110001100101;
		S266reg [LFSR_S-1:0] <= 16'b0100101000010111;
		S267reg [LFSR_S-1:0] <= 16'b0101011010111011;
		S268reg [LFSR_S-1:0] <= 16'b0100000110011011;
		S269reg [LFSR_S-1:0] <= 16'b0000000110100111;
		S270reg [LFSR_S-1:0] <= 16'b0111001010000011;
		S271reg [LFSR_S-1:0] <= 16'b0111111010110100;
		S272reg [LFSR_S-1:0] <= 16'b1010000000000111;
		S273reg [LFSR_S-1:0] <= 16'b0011100111101000;
		S274reg [LFSR_S-1:0] <= 16'b0100110001001000;
		S275reg [LFSR_S-1:0] <= 16'b0111101010111100;
		S276reg [LFSR_S-1:0] <= 16'b0101010110010010;
		S277reg [LFSR_S-1:0] <= 16'b1001101100111000;
		S278reg [LFSR_S-1:0] <= 16'b0000011101110000;
		S279reg [LFSR_S-1:0] <= 16'b1100000110001001;
	end
	if (n1==3) begin
		S0reg [LFSR_S-1:0] <= 16'b0100110000101110;
		S1reg [LFSR_S-1:0] <= 16'b0000101111110110;
		S2reg [LFSR_S-1:0] <= 16'b1111010000101001;
		S3reg [LFSR_S-1:0] <= 16'b0001011101001011;
		S4reg [LFSR_S-1:0] <= 16'b1011001100111111;
		S5reg [LFSR_S-1:0] <= 16'b0001100110001110;
		S6reg [LFSR_S-1:0] <= 16'b1000010111111011;
		S7reg [LFSR_S-1:0] <= 16'b0011001101000100;
		S8reg [LFSR_S-1:0] <= 16'b1110111111010111;
		S9reg [LFSR_S-1:0] <= 16'b0011011101101100;
		S10reg [LFSR_S-1:0] <= 16'b1001111010101101;
		S11reg [LFSR_S-1:0] <= 16'b1110010010100000;
		S12reg [LFSR_S-1:0] <= 16'b1101110100110001;
		S13reg [LFSR_S-1:0] <= 16'b1001001101000111;
		S14reg [LFSR_S-1:0] <= 16'b1111101010000100;
		S15reg [LFSR_S-1:0] <= 16'b1010011000100001;
		S16reg [LFSR_S-1:0] <= 16'b1001011011001101;
		S17reg [LFSR_S-1:0] <= 16'b0110101000100010;
		S18reg [LFSR_S-1:0] <= 16'b0000001011111010;
		S19reg [LFSR_S-1:0] <= 16'b0110110010000011;
		S20reg [LFSR_S-1:0] <= 16'b0001101101111111;
		S21reg [LFSR_S-1:0] <= 16'b1111101010001101;
		S22reg [LFSR_S-1:0] <= 16'b0001001011010010;
		S23reg [LFSR_S-1:0] <= 16'b1111001101001001;
		S24reg [LFSR_S-1:0] <= 16'b0000001000001110;
		S25reg [LFSR_S-1:0] <= 16'b0111011110111010;
		S26reg [LFSR_S-1:0] <= 16'b0011101011111010;
		S27reg [LFSR_S-1:0] <= 16'b0001101011101010;
		S28reg [LFSR_S-1:0] <= 16'b1100010001110101;
		S29reg [LFSR_S-1:0] <= 16'b0011001110100111;
		S30reg [LFSR_S-1:0] <= 16'b1011010011011010;
		S31reg [LFSR_S-1:0] <= 16'b0001110111010011;
		S32reg [LFSR_S-1:0] <= 16'b0011110010000111;
		S33reg [LFSR_S-1:0] <= 16'b1011000110111111;
		S34reg [LFSR_S-1:0] <= 16'b0111010000011001;
		S35reg [LFSR_S-1:0] <= 16'b1001111010110101;
		S36reg [LFSR_S-1:0] <= 16'b0110011111110111;
		S37reg [LFSR_S-1:0] <= 16'b0100010010011100;
		S38reg [LFSR_S-1:0] <= 16'b1010001110000011;
		S39reg [LFSR_S-1:0] <= 16'b0000101101111011;
		S40reg [LFSR_S-1:0] <= 16'b1100100001000101;
		S41reg [LFSR_S-1:0] <= 16'b1110000001101001;
		S42reg [LFSR_S-1:0] <= 16'b0100000010111000;
		S43reg [LFSR_S-1:0] <= 16'b1100101110010011;
		S44reg [LFSR_S-1:0] <= 16'b0101000010111000;
		S45reg [LFSR_S-1:0] <= 16'b1000110011000110;
		S46reg [LFSR_S-1:0] <= 16'b0011001101001110;
		S47reg [LFSR_S-1:0] <= 16'b0100010111110000;
		S48reg [LFSR_S-1:0] <= 16'b1011011100000101;
		S49reg [LFSR_S-1:0] <= 16'b0111011010100110;
		S50reg [LFSR_S-1:0] <= 16'b1101001001000100;
		S51reg [LFSR_S-1:0] <= 16'b0110110111100010;
		S52reg [LFSR_S-1:0] <= 16'b0111101000001000;
		S53reg [LFSR_S-1:0] <= 16'b1011000010001000;
		S54reg [LFSR_S-1:0] <= 16'b1100101111101111;
		S55reg [LFSR_S-1:0] <= 16'b0000110011011111;
		S56reg [LFSR_S-1:0] <= 16'b0011001010100011;
		S57reg [LFSR_S-1:0] <= 16'b0101011100110111;
		S58reg [LFSR_S-1:0] <= 16'b0011001101001100;
		S59reg [LFSR_S-1:0] <= 16'b1100100101100011;
		S60reg [LFSR_S-1:0] <= 16'b0110001001110100;
		S61reg [LFSR_S-1:0] <= 16'b0011101110100010;
		S62reg [LFSR_S-1:0] <= 16'b0001011010101110;
		S63reg [LFSR_S-1:0] <= 16'b1010010111001111;
		S64reg [LFSR_S-1:0] <= 16'b1110011010000100;
		S65reg [LFSR_S-1:0] <= 16'b1101010111111110;
		S66reg [LFSR_S-1:0] <= 16'b1100001111101001;
		S67reg [LFSR_S-1:0] <= 16'b0011001011111010;
		S68reg [LFSR_S-1:0] <= 16'b0000101011111011;
		S69reg [LFSR_S-1:0] <= 16'b0010011101111000;
		S70reg [LFSR_S-1:0] <= 16'b1100011100101111;
		S71reg [LFSR_S-1:0] <= 16'b0100111001111011;
		S72reg [LFSR_S-1:0] <= 16'b0000010001101110;
		S73reg [LFSR_S-1:0] <= 16'b1111001111000011;
		S74reg [LFSR_S-1:0] <= 16'b0101110011001010;
		S75reg [LFSR_S-1:0] <= 16'b1001110010000100;
		S76reg [LFSR_S-1:0] <= 16'b0011001010101001;
		S77reg [LFSR_S-1:0] <= 16'b0110000001001110;
		S78reg [LFSR_S-1:0] <= 16'b1110010111101011;
		S79reg [LFSR_S-1:0] <= 16'b1001101001010111;
		S80reg [LFSR_S-1:0] <= 16'b0101010011111100;
		S81reg [LFSR_S-1:0] <= 16'b1111010010001011;
		S82reg [LFSR_S-1:0] <= 16'b0000100101101010;
		S83reg [LFSR_S-1:0] <= 16'b0111101000111100;
		S84reg [LFSR_S-1:0] <= 16'b1000011100011100;
		S85reg [LFSR_S-1:0] <= 16'b1101111100101011;
		S86reg [LFSR_S-1:0] <= 16'b1011101100001111;
		S87reg [LFSR_S-1:0] <= 16'b0001111010101111;
		S88reg [LFSR_S-1:0] <= 16'b0111001101011000;
		S89reg [LFSR_S-1:0] <= 16'b0000100111111100;
		S90reg [LFSR_S-1:0] <= 16'b0100001011100100;
		S91reg [LFSR_S-1:0] <= 16'b0110001010010010;
		S92reg [LFSR_S-1:0] <= 16'b1001000000000110;
		S93reg [LFSR_S-1:0] <= 16'b1111111110110111;
		S94reg [LFSR_S-1:0] <= 16'b1101000000011010;
		S95reg [LFSR_S-1:0] <= 16'b0111111101001100;
		S96reg [LFSR_S-1:0] <= 16'b0001000001011111;
		S97reg [LFSR_S-1:0] <= 16'b0110000101001011;
		S98reg [LFSR_S-1:0] <= 16'b0011110010111110;
		S99reg [LFSR_S-1:0] <= 16'b1101111101001011;
		S100reg [LFSR_S-1:0] <= 16'b0110000000001000;
		S101reg [LFSR_S-1:0] <= 16'b1110010111000111;
		S102reg [LFSR_S-1:0] <= 16'b1000101100111100;
		S103reg [LFSR_S-1:0] <= 16'b1110001011100101;
		S104reg [LFSR_S-1:0] <= 16'b1110111100011011;
		S105reg [LFSR_S-1:0] <= 16'b1011000101110011;
		S106reg [LFSR_S-1:0] <= 16'b0011100011011110;
		S107reg [LFSR_S-1:0] <= 16'b1000000110110010;
		S108reg [LFSR_S-1:0] <= 16'b0010101011101110;
		S109reg [LFSR_S-1:0] <= 16'b1111010010011111;
		S110reg [LFSR_S-1:0] <= 16'b0111010100000111;
		S111reg [LFSR_S-1:0] <= 16'b0111011111010101;
		S112reg [LFSR_S-1:0] <= 16'b1000110110111011;
		S113reg [LFSR_S-1:0] <= 16'b0011001110101101;
		S114reg [LFSR_S-1:0] <= 16'b0011011111110010;
		S115reg [LFSR_S-1:0] <= 16'b0110111101010010;
		S116reg [LFSR_S-1:0] <= 16'b1101110000101010;
		S117reg [LFSR_S-1:0] <= 16'b0110000001010000;
		S118reg [LFSR_S-1:0] <= 16'b1000010100000010;
		S119reg [LFSR_S-1:0] <= 16'b0110111111000010;
		S120reg [LFSR_S-1:0] <= 16'b1010011011001110;
		S121reg [LFSR_S-1:0] <= 16'b0010101011101001;
		S122reg [LFSR_S-1:0] <= 16'b0001111000100010;
		S123reg [LFSR_S-1:0] <= 16'b1100011100101010;
		S124reg [LFSR_S-1:0] <= 16'b0010000111111100;
		S125reg [LFSR_S-1:0] <= 16'b0111010001101110;
		S126reg [LFSR_S-1:0] <= 16'b1011110000111111;
		S127reg [LFSR_S-1:0] <= 16'b1101101100011011;
		S128reg [LFSR_S-1:0] <= 16'b0100100100101000;
		S129reg [LFSR_S-1:0] <= 16'b1010111101100011;
		S130reg [LFSR_S-1:0] <= 16'b0010111000010010;
		S131reg [LFSR_S-1:0] <= 16'b0110001111100011;
		S132reg [LFSR_S-1:0] <= 16'b0001011101011100;
		S133reg [LFSR_S-1:0] <= 16'b1011011101100101;
		S134reg [LFSR_S-1:0] <= 16'b1001001011000100;
		S135reg [LFSR_S-1:0] <= 16'b0101111101111100;
		S136reg [LFSR_S-1:0] <= 16'b1101010100000111;
		S137reg [LFSR_S-1:0] <= 16'b0100001110001000;
		S138reg [LFSR_S-1:0] <= 16'b0100001001111100;
		S139reg [LFSR_S-1:0] <= 16'b0000111100000101;
	end
	if (n2==3) begin
		S140reg [LFSR_S-1:0] <= 16'b1011100101001101;
		S141reg [LFSR_S-1:0] <= 16'b1010101001101111;
		S142reg [LFSR_S-1:0] <= 16'b1110101011011011;
		S143reg [LFSR_S-1:0] <= 16'b0011001001100010;
		S144reg [LFSR_S-1:0] <= 16'b0101010000011000;
		S145reg [LFSR_S-1:0] <= 16'b0111101110010111;
		S146reg [LFSR_S-1:0] <= 16'b1000110100001100;
		S147reg [LFSR_S-1:0] <= 16'b1110010101100111;
		S148reg [LFSR_S-1:0] <= 16'b0111001011000100;
		S149reg [LFSR_S-1:0] <= 16'b0101000000110110;
		S150reg [LFSR_S-1:0] <= 16'b1001100010000111;
		S151reg [LFSR_S-1:0] <= 16'b0001111101001011;
		S152reg [LFSR_S-1:0] <= 16'b1001110110011111;
		S153reg [LFSR_S-1:0] <= 16'b0000101100101000;
		S154reg [LFSR_S-1:0] <= 16'b1100110111011011;
		S155reg [LFSR_S-1:0] <= 16'b0101001001111000;
		S156reg [LFSR_S-1:0] <= 16'b0111110100110011;
		S157reg [LFSR_S-1:0] <= 16'b1100000010101000;
		S158reg [LFSR_S-1:0] <= 16'b1000100001001111;
		S159reg [LFSR_S-1:0] <= 16'b0111101000100001;
		S160reg [LFSR_S-1:0] <= 16'b1110000001110001;
		S161reg [LFSR_S-1:0] <= 16'b1111110011001011;
		S162reg [LFSR_S-1:0] <= 16'b0111001111010110;
		S163reg [LFSR_S-1:0] <= 16'b1100010111001110;
		S164reg [LFSR_S-1:0] <= 16'b1100000100110000;
		S165reg [LFSR_S-1:0] <= 16'b1111000000101011;
		S166reg [LFSR_S-1:0] <= 16'b0001000010110100;
		S167reg [LFSR_S-1:0] <= 16'b0010000101011111;
		S168reg [LFSR_S-1:0] <= 16'b0011011001000010;
		S169reg [LFSR_S-1:0] <= 16'b1011001111110011;
		S170reg [LFSR_S-1:0] <= 16'b0010111001111101;
		S171reg [LFSR_S-1:0] <= 16'b1010011110110111;
		S172reg [LFSR_S-1:0] <= 16'b0010100101100000;
		S173reg [LFSR_S-1:0] <= 16'b1011101101110001;
		S174reg [LFSR_S-1:0] <= 16'b0111111000010100;
		S175reg [LFSR_S-1:0] <= 16'b0001010111101011;
		S176reg [LFSR_S-1:0] <= 16'b1110110101111101;
		S177reg [LFSR_S-1:0] <= 16'b0001110000000100;
		S178reg [LFSR_S-1:0] <= 16'b1000101110000111;
		S179reg [LFSR_S-1:0] <= 16'b0101001110100100;
		S180reg [LFSR_S-1:0] <= 16'b0010111100011110;
		S181reg [LFSR_S-1:0] <= 16'b0111001010010000;
		S182reg [LFSR_S-1:0] <= 16'b0011011000111000;
		S183reg [LFSR_S-1:0] <= 16'b0111010010110000;
		S184reg [LFSR_S-1:0] <= 16'b1001000110100010;
		S185reg [LFSR_S-1:0] <= 16'b1100111011000100;
		S186reg [LFSR_S-1:0] <= 16'b0101111001101100;
		S187reg [LFSR_S-1:0] <= 16'b0000001100100001;
		S188reg [LFSR_S-1:0] <= 16'b1111111101010111;
		S189reg [LFSR_S-1:0] <= 16'b1000111001000011;
		S190reg [LFSR_S-1:0] <= 16'b1010110100001111;
		S191reg [LFSR_S-1:0] <= 16'b1111101110011011;
		S192reg [LFSR_S-1:0] <= 16'b1100001110100001;
		S193reg [LFSR_S-1:0] <= 16'b1100000110011101;
		S194reg [LFSR_S-1:0] <= 16'b1100011001101100;
		S195reg [LFSR_S-1:0] <= 16'b0000101010110100;
		S196reg [LFSR_S-1:0] <= 16'b0110000101101000;
		S197reg [LFSR_S-1:0] <= 16'b1010000110111010;
		S198reg [LFSR_S-1:0] <= 16'b0000001110000110;
		S199reg [LFSR_S-1:0] <= 16'b0110110011110011;
		S200reg [LFSR_S-1:0] <= 16'b0111111000001001;
		S201reg [LFSR_S-1:0] <= 16'b1111101001100000;
		S202reg [LFSR_S-1:0] <= 16'b1110011110011110;
		S203reg [LFSR_S-1:0] <= 16'b1110011010011000;
		S204reg [LFSR_S-1:0] <= 16'b1111011100010011;
		S205reg [LFSR_S-1:0] <= 16'b0011110010111010;
		S206reg [LFSR_S-1:0] <= 16'b1010001001110110;
		S207reg [LFSR_S-1:0] <= 16'b0000001101101110;
		S208reg [LFSR_S-1:0] <= 16'b1000011110010111;
		S209reg [LFSR_S-1:0] <= 16'b0010100101011000;
		S210reg [LFSR_S-1:0] <= 16'b0011001000100010;
		S211reg [LFSR_S-1:0] <= 16'b1011000011100010;
		S212reg [LFSR_S-1:0] <= 16'b0000110111100000;
		S213reg [LFSR_S-1:0] <= 16'b0000011110100111;
		S214reg [LFSR_S-1:0] <= 16'b0110100111110000;
		S215reg [LFSR_S-1:0] <= 16'b0000010000001110;
		S216reg [LFSR_S-1:0] <= 16'b1010000100010010;
		S217reg [LFSR_S-1:0] <= 16'b1101011010101001;
		S218reg [LFSR_S-1:0] <= 16'b0011110011100101;
		S219reg [LFSR_S-1:0] <= 16'b0000101100001110;
		S220reg [LFSR_S-1:0] <= 16'b0110111010101000;
		S221reg [LFSR_S-1:0] <= 16'b1110001011110001;
		S222reg [LFSR_S-1:0] <= 16'b0010100001010000;
		S223reg [LFSR_S-1:0] <= 16'b1100110111011101;
		S224reg [LFSR_S-1:0] <= 16'b0110011100100010;
		S225reg [LFSR_S-1:0] <= 16'b0110111100100100;
		S226reg [LFSR_S-1:0] <= 16'b0111001100000101;
		S227reg [LFSR_S-1:0] <= 16'b0101100100010011;
		S228reg [LFSR_S-1:0] <= 16'b0010110110101110;
		S229reg [LFSR_S-1:0] <= 16'b1010001110011000;
		S230reg [LFSR_S-1:0] <= 16'b0011010001110010;
		S231reg [LFSR_S-1:0] <= 16'b1111110110001110;
		S232reg [LFSR_S-1:0] <= 16'b0111111101111010;
		S233reg [LFSR_S-1:0] <= 16'b0100101110001000;
		S234reg [LFSR_S-1:0] <= 16'b1000111001000000;
		S235reg [LFSR_S-1:0] <= 16'b1111110111101111;
		S236reg [LFSR_S-1:0] <= 16'b0101010001011011;
		S237reg [LFSR_S-1:0] <= 16'b0100001101110000;
		S238reg [LFSR_S-1:0] <= 16'b0100011100110010;
		S239reg [LFSR_S-1:0] <= 16'b0100011011000110;
		S240reg [LFSR_S-1:0] <= 16'b0001001101001110;
		S241reg [LFSR_S-1:0] <= 16'b1001001010101111;
		S242reg [LFSR_S-1:0] <= 16'b0111000011101101;
		S243reg [LFSR_S-1:0] <= 16'b1000111100100100;
		S244reg [LFSR_S-1:0] <= 16'b0011100101100110;
		S245reg [LFSR_S-1:0] <= 16'b0010001110101010;
		S246reg [LFSR_S-1:0] <= 16'b1000111011101001;
		S247reg [LFSR_S-1:0] <= 16'b0011101101000110;
		S248reg [LFSR_S-1:0] <= 16'b1111110011011100;
		S249reg [LFSR_S-1:0] <= 16'b0111100000110000;
		S250reg [LFSR_S-1:0] <= 16'b0010010111100100;
		S251reg [LFSR_S-1:0] <= 16'b0101011000011010;
		S252reg [LFSR_S-1:0] <= 16'b0010111111101100;
		S253reg [LFSR_S-1:0] <= 16'b0110110000110100;
		S254reg [LFSR_S-1:0] <= 16'b1011101001101111;
		S255reg [LFSR_S-1:0] <= 16'b1000010000101111;
		S256reg [LFSR_S-1:0] <= 16'b1111100100010101;
		S257reg [LFSR_S-1:0] <= 16'b1100011110111001;
		S258reg [LFSR_S-1:0] <= 16'b0011111010111111;
		S259reg [LFSR_S-1:0] <= 16'b0001101010100111;
		S260reg [LFSR_S-1:0] <= 16'b1011100110110001;
		S261reg [LFSR_S-1:0] <= 16'b0101001000010110;
		S262reg [LFSR_S-1:0] <= 16'b0100011100111000;
		S263reg [LFSR_S-1:0] <= 16'b0010101111000010;
		S264reg [LFSR_S-1:0] <= 16'b1001101110010111;
		S265reg [LFSR_S-1:0] <= 16'b1000111111111011;
		S266reg [LFSR_S-1:0] <= 16'b1110000010100010;
		S267reg [LFSR_S-1:0] <= 16'b0000001110100010;
		S268reg [LFSR_S-1:0] <= 16'b1111011011010001;
		S269reg [LFSR_S-1:0] <= 16'b0100011100000000;
		S270reg [LFSR_S-1:0] <= 16'b0000110001101000;
		S271reg [LFSR_S-1:0] <= 16'b0101100100100010;
		S272reg [LFSR_S-1:0] <= 16'b1100011011100011;
		S273reg [LFSR_S-1:0] <= 16'b1010011110110000;
		S274reg [LFSR_S-1:0] <= 16'b1111110100001001;
		S275reg [LFSR_S-1:0] <= 16'b0001101110101000;
		S276reg [LFSR_S-1:0] <= 16'b0011010101000111;
		S277reg [LFSR_S-1:0] <= 16'b1101010000110111;
		S278reg [LFSR_S-1:0] <= 16'b0001001011110001;
		S279reg [LFSR_S-1:0] <= 16'b0110100010101100;
	end
	if (n1==4) begin
		S0reg [LFSR_S-1:0] <= 16'b0100010000000000;
		S1reg [LFSR_S-1:0] <= 16'b0101111101110100;
		S2reg [LFSR_S-1:0] <= 16'b1010100110001000;
		S3reg [LFSR_S-1:0] <= 16'b1001011000001111;
		S4reg [LFSR_S-1:0] <= 16'b0101111010010001;
		S5reg [LFSR_S-1:0] <= 16'b1110101011000001;
		S6reg [LFSR_S-1:0] <= 16'b1111011001011010;
		S7reg [LFSR_S-1:0] <= 16'b1110100111010001;
		S8reg [LFSR_S-1:0] <= 16'b0000100001000001;
		S9reg [LFSR_S-1:0] <= 16'b1001100000110001;
		S10reg [LFSR_S-1:0] <= 16'b0110001111010110;
		S11reg [LFSR_S-1:0] <= 16'b1010001100110101;
		S12reg [LFSR_S-1:0] <= 16'b1101010010001001;
		S13reg [LFSR_S-1:0] <= 16'b0011111110011110;
		S14reg [LFSR_S-1:0] <= 16'b0001001110010010;
		S15reg [LFSR_S-1:0] <= 16'b0100000011110011;
		S16reg [LFSR_S-1:0] <= 16'b0010011111010000;
		S17reg [LFSR_S-1:0] <= 16'b1011101110010000;
		S18reg [LFSR_S-1:0] <= 16'b1111100000010001;
		S19reg [LFSR_S-1:0] <= 16'b0011000010010001;
		S20reg [LFSR_S-1:0] <= 16'b1010000111100010;
		S21reg [LFSR_S-1:0] <= 16'b0001111101011011;
		S22reg [LFSR_S-1:0] <= 16'b1100100000010110;
		S23reg [LFSR_S-1:0] <= 16'b1100010100101001;
		S24reg [LFSR_S-1:0] <= 16'b1110110010101000;
		S25reg [LFSR_S-1:0] <= 16'b1100010011110101;
		S26reg [LFSR_S-1:0] <= 16'b1010000001001011;
		S27reg [LFSR_S-1:0] <= 16'b1001011011100111;
		S28reg [LFSR_S-1:0] <= 16'b1111110111000011;
		S29reg [LFSR_S-1:0] <= 16'b1011101100011011;
		S30reg [LFSR_S-1:0] <= 16'b1100000001111001;
		S31reg [LFSR_S-1:0] <= 16'b1011001000010101;
		S32reg [LFSR_S-1:0] <= 16'b1011111111011001;
		S33reg [LFSR_S-1:0] <= 16'b0101011000111111;
		S34reg [LFSR_S-1:0] <= 16'b1110000110101111;
		S35reg [LFSR_S-1:0] <= 16'b1001000101111001;
		S36reg [LFSR_S-1:0] <= 16'b0111110000101111;
		S37reg [LFSR_S-1:0] <= 16'b1100000010101110;
		S38reg [LFSR_S-1:0] <= 16'b1001010001010000;
		S39reg [LFSR_S-1:0] <= 16'b1001000100010101;
		S40reg [LFSR_S-1:0] <= 16'b0010111000100100;
		S41reg [LFSR_S-1:0] <= 16'b1100001010010000;
		S42reg [LFSR_S-1:0] <= 16'b0000010111111010;
		S43reg [LFSR_S-1:0] <= 16'b0111001000011010;
		S44reg [LFSR_S-1:0] <= 16'b1110101011010011;
		S45reg [LFSR_S-1:0] <= 16'b0101101001111010;
		S46reg [LFSR_S-1:0] <= 16'b0111100101111001;
		S47reg [LFSR_S-1:0] <= 16'b0010010011110000;
		S48reg [LFSR_S-1:0] <= 16'b1111111110111011;
		S49reg [LFSR_S-1:0] <= 16'b0111100010010100;
		S50reg [LFSR_S-1:0] <= 16'b1100010110101001;
		S51reg [LFSR_S-1:0] <= 16'b1111000111100000;
		S52reg [LFSR_S-1:0] <= 16'b1001101110010101;
		S53reg [LFSR_S-1:0] <= 16'b0110110011001010;
		S54reg [LFSR_S-1:0] <= 16'b0001011001001000;
		S55reg [LFSR_S-1:0] <= 16'b1001000011100100;
		S56reg [LFSR_S-1:0] <= 16'b0011100010100111;
		S57reg [LFSR_S-1:0] <= 16'b0001000110000010;
		S58reg [LFSR_S-1:0] <= 16'b0010101100100010;
		S59reg [LFSR_S-1:0] <= 16'b1101100110101100;
		S60reg [LFSR_S-1:0] <= 16'b0101111110001011;
		S61reg [LFSR_S-1:0] <= 16'b0000110101100010;
		S62reg [LFSR_S-1:0] <= 16'b0111000111010010;
		S63reg [LFSR_S-1:0] <= 16'b0100111001010100;
		S64reg [LFSR_S-1:0] <= 16'b0110011111000101;
		S65reg [LFSR_S-1:0] <= 16'b1101100111100110;
		S66reg [LFSR_S-1:0] <= 16'b1000101110101101;
		S67reg [LFSR_S-1:0] <= 16'b1110101011000010;
		S68reg [LFSR_S-1:0] <= 16'b1010111111110001;
		S69reg [LFSR_S-1:0] <= 16'b1011110110101111;
		S70reg [LFSR_S-1:0] <= 16'b0000100010100100;
		S71reg [LFSR_S-1:0] <= 16'b0110100001011101;
		S72reg [LFSR_S-1:0] <= 16'b1110101010001100;
		S73reg [LFSR_S-1:0] <= 16'b1010111011101001;
		S74reg [LFSR_S-1:0] <= 16'b0011110101010010;
		S75reg [LFSR_S-1:0] <= 16'b0000101000101000;
		S76reg [LFSR_S-1:0] <= 16'b0111000000010001;
		S77reg [LFSR_S-1:0] <= 16'b0100111001111000;
		S78reg [LFSR_S-1:0] <= 16'b1001010000000010;
		S79reg [LFSR_S-1:0] <= 16'b1001111011010101;
		S80reg [LFSR_S-1:0] <= 16'b0101111001010000;
		S81reg [LFSR_S-1:0] <= 16'b1101011100000110;
		S82reg [LFSR_S-1:0] <= 16'b0100110000000111;
		S83reg [LFSR_S-1:0] <= 16'b0000100000010100;
		S84reg [LFSR_S-1:0] <= 16'b0100110000011000;
		S85reg [LFSR_S-1:0] <= 16'b0011010100011111;
		S86reg [LFSR_S-1:0] <= 16'b1100111110111011;
		S87reg [LFSR_S-1:0] <= 16'b1111111001100101;
		S88reg [LFSR_S-1:0] <= 16'b0110000011100000;
		S89reg [LFSR_S-1:0] <= 16'b1001111110010101;
		S90reg [LFSR_S-1:0] <= 16'b0101011111111010;
		S91reg [LFSR_S-1:0] <= 16'b0111000110100001;
		S92reg [LFSR_S-1:0] <= 16'b1011011010100111;
		S93reg [LFSR_S-1:0] <= 16'b0100001001100110;
		S94reg [LFSR_S-1:0] <= 16'b1010001111100010;
		S95reg [LFSR_S-1:0] <= 16'b1000011111111101;
		S96reg [LFSR_S-1:0] <= 16'b1111111111010101;
		S97reg [LFSR_S-1:0] <= 16'b0010010001011110;
		S98reg [LFSR_S-1:0] <= 16'b0010000010101010;
		S99reg [LFSR_S-1:0] <= 16'b0010001110011110;
		S100reg [LFSR_S-1:0] <= 16'b0101101000111100;
		S101reg [LFSR_S-1:0] <= 16'b0010011010000000;
		S102reg [LFSR_S-1:0] <= 16'b1010100100110110;
		S103reg [LFSR_S-1:0] <= 16'b0110000000101100;
		S104reg [LFSR_S-1:0] <= 16'b0000100110011011;
		S105reg [LFSR_S-1:0] <= 16'b1101100101010101;
		S106reg [LFSR_S-1:0] <= 16'b1001001010000000;
		S107reg [LFSR_S-1:0] <= 16'b1011000011001111;
		S108reg [LFSR_S-1:0] <= 16'b0000001111000011;
		S109reg [LFSR_S-1:0] <= 16'b1010110000001001;
		S110reg [LFSR_S-1:0] <= 16'b0010010111110001;
		S111reg [LFSR_S-1:0] <= 16'b0101011000001010;
		S112reg [LFSR_S-1:0] <= 16'b1101100001110100;
		S113reg [LFSR_S-1:0] <= 16'b0101001010110001;
		S114reg [LFSR_S-1:0] <= 16'b0101101001101100;
		S115reg [LFSR_S-1:0] <= 16'b0010000101100000;
		S116reg [LFSR_S-1:0] <= 16'b0010100111011010;
		S117reg [LFSR_S-1:0] <= 16'b0001111100011010;
		S118reg [LFSR_S-1:0] <= 16'b1110110101010001;
		S119reg [LFSR_S-1:0] <= 16'b1101000111110101;
		S120reg [LFSR_S-1:0] <= 16'b0001111100000010;
		S121reg [LFSR_S-1:0] <= 16'b1010011001000100;
		S122reg [LFSR_S-1:0] <= 16'b1101101001010111;
		S123reg [LFSR_S-1:0] <= 16'b1111010111111011;
		S124reg [LFSR_S-1:0] <= 16'b1111111111101010;
		S125reg [LFSR_S-1:0] <= 16'b0000011000000010;
		S126reg [LFSR_S-1:0] <= 16'b0111000111010110;
		S127reg [LFSR_S-1:0] <= 16'b0100000110011111;
		S128reg [LFSR_S-1:0] <= 16'b0000111111110101;
		S129reg [LFSR_S-1:0] <= 16'b0111010001101111;
		S130reg [LFSR_S-1:0] <= 16'b1000011101000100;
		S131reg [LFSR_S-1:0] <= 16'b1011011011001101;
		S132reg [LFSR_S-1:0] <= 16'b0111000001110110;
		S133reg [LFSR_S-1:0] <= 16'b1000100110010000;
		S134reg [LFSR_S-1:0] <= 16'b0011010110000010;
		S135reg [LFSR_S-1:0] <= 16'b1010101001011101;
		S136reg [LFSR_S-1:0] <= 16'b1101110100011111;
		S137reg [LFSR_S-1:0] <= 16'b1111010111010000;
		S138reg [LFSR_S-1:0] <= 16'b0111101101010010;
		S139reg [LFSR_S-1:0] <= 16'b0100001101101000;
	end
	if (n2==4) begin
		S140reg [LFSR_S-1:0] <= 16'b1110100111100101;
		S141reg [LFSR_S-1:0] <= 16'b1001110011000111;
		S142reg [LFSR_S-1:0] <= 16'b1101111000001011;
		S143reg [LFSR_S-1:0] <= 16'b0100001111010110;
		S144reg [LFSR_S-1:0] <= 16'b0111011010100110;
		S145reg [LFSR_S-1:0] <= 16'b0001100111110110;
		S146reg [LFSR_S-1:0] <= 16'b1111000111001101;
		S147reg [LFSR_S-1:0] <= 16'b0011100011100010;
		S148reg [LFSR_S-1:0] <= 16'b1100011111100011;
		S149reg [LFSR_S-1:0] <= 16'b1101001011000011;
		S150reg [LFSR_S-1:0] <= 16'b1001010111010110;
		S151reg [LFSR_S-1:0] <= 16'b0010001111111101;
		S152reg [LFSR_S-1:0] <= 16'b0100110110010100;
		S153reg [LFSR_S-1:0] <= 16'b1110110100111101;
		S154reg [LFSR_S-1:0] <= 16'b0010101101000110;
		S155reg [LFSR_S-1:0] <= 16'b1100100100000100;
		S156reg [LFSR_S-1:0] <= 16'b0111111010001110;
		S157reg [LFSR_S-1:0] <= 16'b0000010100011100;
		S158reg [LFSR_S-1:0] <= 16'b0010100110101110;
		S159reg [LFSR_S-1:0] <= 16'b1101111110010000;
		S160reg [LFSR_S-1:0] <= 16'b1100010100001111;
		S161reg [LFSR_S-1:0] <= 16'b1001000010101001;
		S162reg [LFSR_S-1:0] <= 16'b0001010100011100;
		S163reg [LFSR_S-1:0] <= 16'b1010010011101010;
		S164reg [LFSR_S-1:0] <= 16'b1011100011111011;
		S165reg [LFSR_S-1:0] <= 16'b0011010000111000;
		S166reg [LFSR_S-1:0] <= 16'b0110111010100100;
		S167reg [LFSR_S-1:0] <= 16'b0101010010010110;
		S168reg [LFSR_S-1:0] <= 16'b0111101100111101;
		S169reg [LFSR_S-1:0] <= 16'b0001100001111001;
		S170reg [LFSR_S-1:0] <= 16'b1011001110101001;
		S171reg [LFSR_S-1:0] <= 16'b0011000011100000;
		S172reg [LFSR_S-1:0] <= 16'b1100001001111101;
		S173reg [LFSR_S-1:0] <= 16'b1100110100010111;
		S174reg [LFSR_S-1:0] <= 16'b1011001000010110;
		S175reg [LFSR_S-1:0] <= 16'b1001100010111100;
		S176reg [LFSR_S-1:0] <= 16'b0110100000101010;
		S177reg [LFSR_S-1:0] <= 16'b0100001101111100;
		S178reg [LFSR_S-1:0] <= 16'b1011001000001001;
		S179reg [LFSR_S-1:0] <= 16'b0101111101110111;
		S180reg [LFSR_S-1:0] <= 16'b1101010101111011;
		S181reg [LFSR_S-1:0] <= 16'b0100000010000101;
		S182reg [LFSR_S-1:0] <= 16'b0101110101111011;
		S183reg [LFSR_S-1:0] <= 16'b0111111110101111;
		S184reg [LFSR_S-1:0] <= 16'b0011111000111001;
		S185reg [LFSR_S-1:0] <= 16'b0001100101110110;
		S186reg [LFSR_S-1:0] <= 16'b1000001010111111;
		S187reg [LFSR_S-1:0] <= 16'b1000111101011111;
		S188reg [LFSR_S-1:0] <= 16'b1111001100010101;
		S189reg [LFSR_S-1:0] <= 16'b0100111011111010;
		S190reg [LFSR_S-1:0] <= 16'b0111010110001100;
		S191reg [LFSR_S-1:0] <= 16'b1100001101100011;
		S192reg [LFSR_S-1:0] <= 16'b0010010101101101;
		S193reg [LFSR_S-1:0] <= 16'b0000111101110011;
		S194reg [LFSR_S-1:0] <= 16'b1010001101100100;
		S195reg [LFSR_S-1:0] <= 16'b1101000001000001;
		S196reg [LFSR_S-1:0] <= 16'b1101101001010011;
		S197reg [LFSR_S-1:0] <= 16'b1010101001111111;
		S198reg [LFSR_S-1:0] <= 16'b0110101011111010;
		S199reg [LFSR_S-1:0] <= 16'b0010001001111010;
		S200reg [LFSR_S-1:0] <= 16'b0101011010011101;
		S201reg [LFSR_S-1:0] <= 16'b1100011101111111;
		S202reg [LFSR_S-1:0] <= 16'b1001111010101111;
		S203reg [LFSR_S-1:0] <= 16'b1011110101011110;
		S204reg [LFSR_S-1:0] <= 16'b1110001110110011;
		S205reg [LFSR_S-1:0] <= 16'b1111011001011010;
		S206reg [LFSR_S-1:0] <= 16'b0101100100000110;
		S207reg [LFSR_S-1:0] <= 16'b1100101100111101;
		S208reg [LFSR_S-1:0] <= 16'b1010011111100100;
		S209reg [LFSR_S-1:0] <= 16'b1101010100000010;
		S210reg [LFSR_S-1:0] <= 16'b0000010011110000;
		S211reg [LFSR_S-1:0] <= 16'b1101111101011011;
		S212reg [LFSR_S-1:0] <= 16'b0010001101000001;
		S213reg [LFSR_S-1:0] <= 16'b1100100111100010;
		S214reg [LFSR_S-1:0] <= 16'b1101101001000010;
		S215reg [LFSR_S-1:0] <= 16'b1001101011011100;
		S216reg [LFSR_S-1:0] <= 16'b1010101101110010;
		S217reg [LFSR_S-1:0] <= 16'b0011110010101111;
		S218reg [LFSR_S-1:0] <= 16'b1110010100111101;
		S219reg [LFSR_S-1:0] <= 16'b1010001101000100;
		S220reg [LFSR_S-1:0] <= 16'b1111000011000101;
		S221reg [LFSR_S-1:0] <= 16'b0100001110101000;
		S222reg [LFSR_S-1:0] <= 16'b1011001100111111;
		S223reg [LFSR_S-1:0] <= 16'b0011111100101110;
		S224reg [LFSR_S-1:0] <= 16'b0110111001111010;
		S225reg [LFSR_S-1:0] <= 16'b1001111110001011;
		S226reg [LFSR_S-1:0] <= 16'b1010101000000001;
		S227reg [LFSR_S-1:0] <= 16'b0001000100011100;
		S228reg [LFSR_S-1:0] <= 16'b0101110010010110;
		S229reg [LFSR_S-1:0] <= 16'b1011111110101001;
		S230reg [LFSR_S-1:0] <= 16'b0010010011001000;
		S231reg [LFSR_S-1:0] <= 16'b0101111110010000;
		S232reg [LFSR_S-1:0] <= 16'b0110101110100010;
		S233reg [LFSR_S-1:0] <= 16'b0000101111011101;
		S234reg [LFSR_S-1:0] <= 16'b1010100011010010;
		S235reg [LFSR_S-1:0] <= 16'b0101101101010101;
		S236reg [LFSR_S-1:0] <= 16'b1001001110110011;
		S237reg [LFSR_S-1:0] <= 16'b0111001010100111;
		S238reg [LFSR_S-1:0] <= 16'b1001111101101101;
		S239reg [LFSR_S-1:0] <= 16'b1000011100000001;
		S240reg [LFSR_S-1:0] <= 16'b0110101101001111;
		S241reg [LFSR_S-1:0] <= 16'b1000010101001011;
		S242reg [LFSR_S-1:0] <= 16'b0111000101110110;
		S243reg [LFSR_S-1:0] <= 16'b1000000011011100;
		S244reg [LFSR_S-1:0] <= 16'b1101011000111101;
		S245reg [LFSR_S-1:0] <= 16'b0001110110110110;
		S246reg [LFSR_S-1:0] <= 16'b1000010011111011;
		S247reg [LFSR_S-1:0] <= 16'b1001110110110110;
		S248reg [LFSR_S-1:0] <= 16'b1100011111010111;
		S249reg [LFSR_S-1:0] <= 16'b0011100010100000;
		S250reg [LFSR_S-1:0] <= 16'b0001111101001110;
		S251reg [LFSR_S-1:0] <= 16'b0010111011110010;
		S252reg [LFSR_S-1:0] <= 16'b0101010010110010;
		S253reg [LFSR_S-1:0] <= 16'b1011011110100011;
		S254reg [LFSR_S-1:0] <= 16'b0110111110001000;
		S255reg [LFSR_S-1:0] <= 16'b0010001001100011;
		S256reg [LFSR_S-1:0] <= 16'b1001110110001101;
		S257reg [LFSR_S-1:0] <= 16'b0001001010111011;
		S258reg [LFSR_S-1:0] <= 16'b0110011110001100;
		S259reg [LFSR_S-1:0] <= 16'b0101100101011011;
		S260reg [LFSR_S-1:0] <= 16'b1100000000110110;
		S261reg [LFSR_S-1:0] <= 16'b1010100110100011;
		S262reg [LFSR_S-1:0] <= 16'b0000011111101110;
		S263reg [LFSR_S-1:0] <= 16'b0001111110011011;
		S264reg [LFSR_S-1:0] <= 16'b0111111011110000;
		S265reg [LFSR_S-1:0] <= 16'b0011000111100100;
		S266reg [LFSR_S-1:0] <= 16'b0011110011000010;
		S267reg [LFSR_S-1:0] <= 16'b1101011110001101;
		S268reg [LFSR_S-1:0] <= 16'b0101010100100110;
		S269reg [LFSR_S-1:0] <= 16'b0010111001100100;
		S270reg [LFSR_S-1:0] <= 16'b0000100010000000;
		S271reg [LFSR_S-1:0] <= 16'b1111001101011101;
		S272reg [LFSR_S-1:0] <= 16'b1101011011110111;
		S273reg [LFSR_S-1:0] <= 16'b0100011101000010;
		S274reg [LFSR_S-1:0] <= 16'b1101010101001000;
		S275reg [LFSR_S-1:0] <= 16'b0111111101001100;
		S276reg [LFSR_S-1:0] <= 16'b0110011101101011;
		S277reg [LFSR_S-1:0] <= 16'b1110001100101100;
		S278reg [LFSR_S-1:0] <= 16'b1111011101011010;
		S279reg [LFSR_S-1:0] <= 16'b1011011100100011;
	end
end
endmodule