// Chris Ceroici

// Stochastic bit generators 

module STOCH(
	PD0, PD1, PD2, PD3, PD4, PD5, PD6, PD7, PD8, PD9, PD10, PD11, PD12, PD13, PD14, PD15, PD16, PD17, PD18, PD19, PD20, PD21, PD22, PD23, PD24, PD25, PD26, PD27, PD28, PD29, PD30, PD31, PD32, PD33, PD34, PD35, PD36, PD37, PD38, PD39, PD40, PD41, PD42, PD43, PD44, PD45, PD46, PD47, PD48, PD49, PD50, PD51, PD52, PD53, PD54, PD55, PD56, PD57, PD58, PD59, PD60, PD61, PD62, PD63, PD64, PD65, PD66, PD67, PD68, PD69, PD70, PD71, PD72, PD73, PD74, PD75, PD76, PD77, PD78, PD79, PD80, PD81, PD82, PD83, PD84, PD85, PD86, PD87, PD88, PD89, PD90, PD91, PD92, PD93, PD94, PD95, PD96, PD97, PD98, PD99, PD100, PD101, PD102, PD103, PD104, PD105, PD106, PD107, PD108, PD109, PD110, PD111, PD112, PD113, PD114, PD115, PD116, PD117, PD118, PD119, PD120, PD121, PD122, PD123, PD124, PD125, PD126, PD127, PD128, PD129, PD130, PD131, PD132, PD133, PD134, PD135, PD136, PD137, PD138, PD139, PD140, PD141, PD142, PD143, PD144, PD145, PD146, PD147, PD148, PD149, PD150, PD151, PD152, PD153, PD154, PD155, PD156, PD157, PD158, PD159, PD160, PD161, PD162, PD163, PD164, PD165, PD166, PD167, PD168, PD169, PD170, PD171, PD172, PD173, PD174, PD175, PD176, PD177, PD178, PD179, PD180, PD181, PD182, PD183, PD184, PD185, PD186, PD187, PD188, PD189, PD190, PD191, PD192, PD193, PD194, PD195, PD196, PD197, PD198, PD199, PD200, PD201, PD202, PD203, PD204, PD205, PD206, PD207, PD208, PD209, PD210, PD211, PD212, PD213, PD214, PD215, PD216, PD217, PD218, PD219, PD220, PD221, PD222, PD223, PD224, PD225, PD226, PD227, PD228, PD229, PD230, PD231, PD232, PD233, PD234, PD235, PD236, PD237, PD238, PD239, PD240, PD241, PD242, PD243, PD244, PD245, PD246, PD247, PD248, PD249, PD250, PD251, PD252, PD253, PD254, PD255, PD256, PD257, PD258, PD259, PD260, PD261, PD262, PD263, PD264, PD265, PD266, PD267, PD268, PD269, PD270, PD271, PD272, PD273, PD274, PD275, PD276, PD277, PD278, PD279, PD280, PD281, PD282, PD283, PD284, PD285, PD286, PD287, PD288, PD289, PD290, PD291, PD292, PD293, PD294, PD295, PD296, PD297, PD298, PD299, PD300, PD301, PD302, PD303, PD304, PD305, PD306, PD307, PD308, PD309, PD310, PD311, PD312, PD313, PD314, PD315, PD316, PD317, PD318, PD319, PD320, PD321, PD322, PD323, PD324, PD325, PD326, PD327, PD328, PD329, PD330, PD331, PD332, PD333, PD334, PD335, PD336, PD337, PD338, PD339, PD340, PD341, PD342, PD343, PD344, PD345, PD346, PD347, PD348, PD349, PD350, PD351, PD352, PD353, PD354, PD355, PD356, PD357, PD358, PD359, PD360, PD361, PD362, PD363, PD364, PD365, PD366, PD367, PD368, PD369, PD370, PD371, PD372, PD373, PD374, PD375, PD376, PD377, PD378, PD379, PD380, PD381, PD382, PD383, PD384, PD385, PD386, PD387, PD388, PD389, PD390, PD391, PD392, PD393, PD394, PD395, PD396, PD397, PD398, PD399, PD400, PD401, PD402, PD403, PD404, PD405, PD406, PD407, PD408, PD409, PD410, PD411, PD412, PD413, PD414, PD415, PD416, PD417, PD418, PD419, PD420, PD421, PD422, PD423, PD424, PD425, PD426, PD427, PD428, PD429, PD430, PD431, PD432, PD433, PD434, PD435, PD436, PD437, PD438, PD439, PD440, PD441, PD442, PD443, PD444, PD445, PD446, PD447, PD448, PD449, PD450, PD451, PD452, PD453, PD454, PD455, PD456,
	PD_long0, PD_long1, PD_long2, PD_long3, PD_long4, PD_long5, PD_long6, PD_long7, PD_long8, PD_long9, PD_long10, PD_long11, PD_long12, PD_long13, PD_long14,
	R0, R1, R2, R3, R4, R5, R6, R7, R8, R9, R10, R11, R12, R13, R14, R15, R16, R17, R18, R19, R20, R21, R22, R23, R24, R25, R26, R27, R28, R29, R30, R31, R32, R33, R34, R35, R36, R37, R38, R39, R40, R41, R42, R43, R44, R45, R46, R47, R48, R49, R50, R51, R52, R53, R54, R55, R56, R57, R58, R59, R60, R61, R62, R63, R64, R65, R66, R67, R68, R69, R70, R71, R72, R73, R74, R75, R76, R77, R78, R79, R80, R81, R82, R83, R84, R85, R86, R87, R88, R89, R90, R91, R92, R93, R94, R95, R96, R97, R98, R99, R100, R101, R102, R103, R104, R105, R106, R107, R108, R109, R110, R111, R112, R113, R114, R115, R116, R117, R118, R119, R120, R121, R122, R123, R124, R125, R126, R127, R128, R129, R130, R131, R132, R133, R134, R135, R136, R137, R138, R139, R140, R141, R142, R143, R144, R145, R146, R147, R148, R149, R150, R151, R152, R153, R154, R155, R156, R157, R158, R159, R160, R161, R162, R163, R164, R165, R166, R167, R168, R169, R170, R171, R172, R173, R174, R175, R176, R177, R178, R179, R180, R181, R182, R183, R184, R185, R186, R187, R188, R189, R190, R191, R192, R193, R194, R195, R196, R197, R198, R199, R200, R201, R202, R203, R204, R205, R206, R207, R208, R209, R210, R211, R212, R213, R214, R215, R216, R217, R218, R219, R220, R221, R222, R223, R224, R225, R226, R227, R228, R229, R230, R231, R232, R233, R234, R235, R236, R237, R238, R239, R240, R241, R242, R243, R244, R245, R246, R247, R248, R249, R250, R251, R252, R253, R254, R255, R256, R257, R258, R259, R260, R261, R262, R263, R264, R265, R266, R267, R268, R269, R270, R271, R272, R273, R274, R275, R276, R277, R278, R279, R280, R281, R282, R283, R284, R285, R286, R287, R288, R289, R290, R291, R292, R293, R294, R295, R296, R297, R298, R299, R300, R301, R302, R303, R304, R305, R306, R307, R308, R309, R310, R311, R312, R313, R314, R315, R316, R317, R318, R319, R320, R321, R322, R323, R324, R325, R326, R327, R328, R329, R330, R331, R332, R333, R334, R335, R336, R337, R338, R339, R340, R341, R342, R343, R344, R345, R346, R347, R348, R349, R350, R351, R352, R353, R354, R355, R356, R357, R358, R359, R360, R361, R362, R363, R364, R365, R366, R367, R368, R369, R370, R371, R372, R373, R374, R375, R376, R377, R378, R379, R380, R381, R382, R383, R384, R385, R386, R387, R388, R389, R390, R391, R392, R393, R394, R395, R396, R397, R398, R399, R400, R401, R402, R403, R404, R405, R406, R407, R408, R409, R410, R411, R412, R413, R414, R415, R416, R417, R418, R419, R420, R421, R422, R423, R424, R425, R426, R427, R428, R429, R430, R431, R432, R433, R434, R435, R436, R437, R438, R439, R440, R441, R442, R443, R444, R445, R446, R447, R448, R449, R450, R451, R452, R453, R454, R455, R456,
	R_long0, R_long1, R_long2, R_long3, R_long4, R_long5, R_long6, R_long7, R_long8, R_long9, R_long10, R_long11, R_long12, R_long13, R_long14,
	P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, P52, P53, P54, P55, P56, P57, P58, P59, P60, P61, P62, P63, P64, P65, P66, P67, P68, P69, P70, P71, P72, P73, P74, P75, P76, P77, P78, P79, P80, P81, P82, P83, P84, P85, P86, P87, P88, P89, P90, P91, P92, P93, P94, P95, P96, P97, P98, P99, P100, P101, P102, P103, P104, P105, P106, P107, P108, P109, P110, P111, P112, P113, P114, P115, P116, P117, P118, P119, P120, P121, P122, P123, P124, P125, P126, P127, P128, P129, P130, P131, P132, P133, P134, P135, P136, P137, P138, P139, P140, P141, P142, P143, P144, P145, P146, P147, P148, P149, P150, P151, P152, P153, P154, P155, P156, P157, P158, P159, P160, P161, P162, P163, P164, P165, P166, P167, P168, P169, P170, P171, P172, P173, P174, P175, P176, P177, P178, P179, P180, P181, P182, P183, P184, P185, P186, P187, P188, P189, P190, P191, P192, P193, P194, P195, P196, P197, P198, P199, P200, P201, P202, P203, P204, P205, P206, P207, P208, P209, P210, P211, P212, P213, P214, P215, P216, P217, P218, P219, P220, P221, P222, P223, P224, P225, P226, P227, P228, P229, P230, P231, P232, P233, P234, P235, P236, P237, P238, P239, P240, P241, P242, P243, P244, P245, P246, P247, P248, P249, P250, P251, P252, P253, P254, P255, P256, P257, P258, P259, P260, P261, P262, P263, P264, P265, P266, P267, P268, P269, P270, P271, P272, P273, P274, P275, P276, P277, P278, P279, P280, P281, P282, P283, P284, P285, P286, P287, P288, P289, P290, P291, P292, P293, P294, P295, P296, P297, P298, P299, P300, P301, P302, P303, P304, P305, P306, P307, P308, P309, P310, P311, P312, P313, P314, P315, P316, P317, P318, P319, P320, P321, P322, P323, P324, P325, P326, P327, P328, P329, P330, P331, P332, P333, P334, P335, P336, P337, P338, P339, P340, P341, P342, P343, P344, P345, P346, P347, P348, P349, P350, P351, P352, P353, P354, P355, P356, P357, P358, P359, P360, P361, P362, P363, P364, P365, P366, P367, P368, P369, P370, P371, P372, P373, P374, P375, P376, P377, P378, P379, P380, P381, P382, P383, P384, P385, P386, P387, P388, P389, P390, P391, P392, P393, P394, P395, P396, P397, P398, P399, P400, P401, P402, P403, P404, P405, P406, P407, P408, P409, P410, P411, P412, P413, P414, P415, P416, P417, P418, P419, P420, P421, P422, P423, P424, P425, P426, P427, P428, P429, P430, P431, P432, P433, P434, P435, P436, P437, P438, P439, P440, P441, P442, P443, P444, P445, P446, P447, P448, P449, P450, P451, P452, P453, P454, P455, P456,
	P_long0, P_long1, P_long2, P_long3, P_long4, P_long5, P_long6, P_long7, P_long8, P_long9, P_long10, P_long11, P_long12, P_long13, P_long14,
	CLK
);

parameter DP_in = 8; // Short Decimal precision 

parameter DP_out = 16; // Long Decimal precision 

input CLK; // Trigger
input wire [DP_in - 1:0] PD0, PD1, PD2, PD3, PD4, PD5, PD6, PD7, PD8, PD9, PD10, PD11, PD12, PD13, PD14, PD15, PD16, PD17, PD18, PD19, PD20, PD21, PD22, PD23, PD24, PD25, PD26, PD27, PD28, PD29, PD30, PD31, PD32, PD33, PD34, PD35, PD36, PD37, PD38, PD39, PD40, PD41, PD42, PD43, PD44, PD45, PD46, PD47, PD48, PD49, PD50, PD51, PD52, PD53, PD54, PD55, PD56, PD57, PD58, PD59, PD60, PD61, PD62, PD63, PD64, PD65, PD66, PD67, PD68, PD69, PD70, PD71, PD72, PD73, PD74, PD75, PD76, PD77, PD78, PD79, PD80, PD81, PD82, PD83, PD84, PD85, PD86, PD87, PD88, PD89, PD90, PD91, PD92, PD93, PD94, PD95, PD96, PD97, PD98, PD99, PD100, PD101, PD102, PD103, PD104, PD105, PD106, PD107, PD108, PD109, PD110, PD111, PD112, PD113, PD114, PD115, PD116, PD117, PD118, PD119, PD120, PD121, PD122, PD123, PD124, PD125, PD126, PD127, PD128, PD129, PD130, PD131, PD132, PD133, PD134, PD135, PD136, PD137, PD138, PD139, PD140, PD141, PD142, PD143, PD144, PD145, PD146, PD147, PD148, PD149, PD150, PD151, PD152, PD153, PD154, PD155, PD156, PD157, PD158, PD159, PD160, PD161, PD162, PD163, PD164, PD165, PD166, PD167, PD168, PD169, PD170, PD171, PD172, PD173, PD174, PD175, PD176, PD177, PD178, PD179, PD180, PD181, PD182, PD183, PD184, PD185, PD186, PD187, PD188, PD189, PD190, PD191, PD192, PD193, PD194, PD195, PD196, PD197, PD198, PD199, PD200, PD201, PD202, PD203, PD204, PD205, PD206, PD207, PD208, PD209, PD210, PD211, PD212, PD213, PD214, PD215, PD216, PD217, PD218, PD219, PD220, PD221, PD222, PD223, PD224, PD225, PD226, PD227, PD228, PD229, PD230, PD231, PD232, PD233, PD234, PD235, PD236, PD237, PD238, PD239, PD240, PD241, PD242, PD243, PD244, PD245, PD246, PD247, PD248, PD249, PD250, PD251, PD252, PD253, PD254, PD255, PD256, PD257, PD258, PD259, PD260, PD261, PD262, PD263, PD264, PD265, PD266, PD267, PD268, PD269, PD270, PD271, PD272, PD273, PD274, PD275, PD276, PD277, PD278, PD279, PD280, PD281, PD282, PD283, PD284, PD285, PD286, PD287, PD288, PD289, PD290, PD291, PD292, PD293, PD294, PD295, PD296, PD297, PD298, PD299, PD300, PD301, PD302, PD303, PD304, PD305, PD306, PD307, PD308, PD309, PD310, PD311, PD312, PD313, PD314, PD315, PD316, PD317, PD318, PD319, PD320, PD321, PD322, PD323, PD324, PD325, PD326, PD327, PD328, PD329, PD330, PD331, PD332, PD333, PD334, PD335, PD336, PD337, PD338, PD339, PD340, PD341, PD342, PD343, PD344, PD345, PD346, PD347, PD348, PD349, PD350, PD351, PD352, PD353, PD354, PD355, PD356, PD357, PD358, PD359, PD360, PD361, PD362, PD363, PD364, PD365, PD366, PD367, PD368, PD369, PD370, PD371, PD372, PD373, PD374, PD375, PD376, PD377, PD378, PD379, PD380, PD381, PD382, PD383, PD384, PD385, PD386, PD387, PD388, PD389, PD390, PD391, PD392, PD393, PD394, PD395, PD396, PD397, PD398, PD399, PD400, PD401, PD402, PD403, PD404, PD405, PD406, PD407, PD408, PD409, PD410, PD411, PD412, PD413, PD414, PD415, PD416, PD417, PD418, PD419, PD420, PD421, PD422, PD423, PD424, PD425, PD426, PD427, PD428, PD429, PD430, PD431, PD432, PD433, PD434, PD435, PD436, PD437, PD438, PD439, PD440, PD441, PD442, PD443, PD444, PD445, PD446, PD447, PD448, PD449, PD450, PD451, PD452, PD453, PD454, PD455, PD456;
input wire [DP_out - 1:0] PD_long0, PD_long1, PD_long2, PD_long3, PD_long4, PD_long5, PD_long6, PD_long7, PD_long8, PD_long9, PD_long10, PD_long11, PD_long12, PD_long13, PD_long14;
input wire [DP_in - 1:0] R0, R1, R2, R3, R4, R5, R6, R7, R8, R9, R10, R11, R12, R13, R14, R15, R16, R17, R18, R19, R20, R21, R22, R23, R24, R25, R26, R27, R28, R29, R30, R31, R32, R33, R34, R35, R36, R37, R38, R39, R40, R41, R42, R43, R44, R45, R46, R47, R48, R49, R50, R51, R52, R53, R54, R55, R56, R57, R58, R59, R60, R61, R62, R63, R64, R65, R66, R67, R68, R69, R70, R71, R72, R73, R74, R75, R76, R77, R78, R79, R80, R81, R82, R83, R84, R85, R86, R87, R88, R89, R90, R91, R92, R93, R94, R95, R96, R97, R98, R99, R100, R101, R102, R103, R104, R105, R106, R107, R108, R109, R110, R111, R112, R113, R114, R115, R116, R117, R118, R119, R120, R121, R122, R123, R124, R125, R126, R127, R128, R129, R130, R131, R132, R133, R134, R135, R136, R137, R138, R139, R140, R141, R142, R143, R144, R145, R146, R147, R148, R149, R150, R151, R152, R153, R154, R155, R156, R157, R158, R159, R160, R161, R162, R163, R164, R165, R166, R167, R168, R169, R170, R171, R172, R173, R174, R175, R176, R177, R178, R179, R180, R181, R182, R183, R184, R185, R186, R187, R188, R189, R190, R191, R192, R193, R194, R195, R196, R197, R198, R199, R200, R201, R202, R203, R204, R205, R206, R207, R208, R209, R210, R211, R212, R213, R214, R215, R216, R217, R218, R219, R220, R221, R222, R223, R224, R225, R226, R227, R228, R229, R230, R231, R232, R233, R234, R235, R236, R237, R238, R239, R240, R241, R242, R243, R244, R245, R246, R247, R248, R249, R250, R251, R252, R253, R254, R255, R256, R257, R258, R259, R260, R261, R262, R263, R264, R265, R266, R267, R268, R269, R270, R271, R272, R273, R274, R275, R276, R277, R278, R279, R280, R281, R282, R283, R284, R285, R286, R287, R288, R289, R290, R291, R292, R293, R294, R295, R296, R297, R298, R299, R300, R301, R302, R303, R304, R305, R306, R307, R308, R309, R310, R311, R312, R313, R314, R315, R316, R317, R318, R319, R320, R321, R322, R323, R324, R325, R326, R327, R328, R329, R330, R331, R332, R333, R334, R335, R336, R337, R338, R339, R340, R341, R342, R343, R344, R345, R346, R347, R348, R349, R350, R351, R352, R353, R354, R355, R356, R357, R358, R359, R360, R361, R362, R363, R364, R365, R366, R367, R368, R369, R370, R371, R372, R373, R374, R375, R376, R377, R378, R379, R380, R381, R382, R383, R384, R385, R386, R387, R388, R389, R390, R391, R392, R393, R394, R395, R396, R397, R398, R399, R400, R401, R402, R403, R404, R405, R406, R407, R408, R409, R410, R411, R412, R413, R414, R415, R416, R417, R418, R419, R420, R421, R422, R423, R424, R425, R426, R427, R428, R429, R430, R431, R432, R433, R434, R435, R436, R437, R438, R439, R440, R441, R442, R443, R444, R445, R446, R447, R448, R449, R450, R451, R452, R453, R454, R455, R456;
input wire [DP_out - 1:0] R_long0, R_long1, R_long2, R_long3, R_long4, R_long5, R_long6, R_long7, R_long8, R_long9, R_long10, R_long11, R_long12, R_long13, R_long14;

output wire P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, P31, P32, P33, P34, P35, P36, P37, P38, P39, P40, P41, P42, P43, P44, P45, P46, P47, P48, P49, P50, P51, P52, P53, P54, P55, P56, P57, P58, P59, P60, P61, P62, P63, P64, P65, P66, P67, P68, P69, P70, P71, P72, P73, P74, P75, P76, P77, P78, P79, P80, P81, P82, P83, P84, P85, P86, P87, P88, P89, P90, P91, P92, P93, P94, P95, P96, P97, P98, P99, P100, P101, P102, P103, P104, P105, P106, P107, P108, P109, P110, P111, P112, P113, P114, P115, P116, P117, P118, P119, P120, P121, P122, P123, P124, P125, P126, P127, P128, P129, P130, P131, P132, P133, P134, P135, P136, P137, P138, P139, P140, P141, P142, P143, P144, P145, P146, P147, P148, P149, P150, P151, P152, P153, P154, P155, P156, P157, P158, P159, P160, P161, P162, P163, P164, P165, P166, P167, P168, P169, P170, P171, P172, P173, P174, P175, P176, P177, P178, P179, P180, P181, P182, P183, P184, P185, P186, P187, P188, P189, P190, P191, P192, P193, P194, P195, P196, P197, P198, P199, P200, P201, P202, P203, P204, P205, P206, P207, P208, P209, P210, P211, P212, P213, P214, P215, P216, P217, P218, P219, P220, P221, P222, P223, P224, P225, P226, P227, P228, P229, P230, P231, P232, P233, P234, P235, P236, P237, P238, P239, P240, P241, P242, P243, P244, P245, P246, P247, P248, P249, P250, P251, P252, P253, P254, P255, P256, P257, P258, P259, P260, P261, P262, P263, P264, P265, P266, P267, P268, P269, P270, P271, P272, P273, P274, P275, P276, P277, P278, P279, P280, P281, P282, P283, P284, P285, P286, P287, P288, P289, P290, P291, P292, P293, P294, P295, P296, P297, P298, P299, P300, P301, P302, P303, P304, P305, P306, P307, P308, P309, P310, P311, P312, P313, P314, P315, P316, P317, P318, P319, P320, P321, P322, P323, P324, P325, P326, P327, P328, P329, P330, P331, P332, P333, P334, P335, P336, P337, P338, P339, P340, P341, P342, P343, P344, P345, P346, P347, P348, P349, P350, P351, P352, P353, P354, P355, P356, P357, P358, P359, P360, P361, P362, P363, P364, P365, P366, P367, P368, P369, P370, P371, P372, P373, P374, P375, P376, P377, P378, P379, P380, P381, P382, P383, P384, P385, P386, P387, P388, P389, P390, P391, P392, P393, P394, P395, P396, P397, P398, P399, P400, P401, P402, P403, P404, P405, P406, P407, P408, P409, P410, P411, P412, P413, P414, P415, P416, P417, P418, P419, P420, P421, P422, P423, P424, P425, P426, P427, P428, P429, P430, P431, P432, P433, P434, P435, P436, P437, P438, P439, P440, P441, P442, P443, P444, P445, P446, P447, P448, P449, P450, P451, P452, P453, P454, P455, P456;
output wire P_long0, P_long1, P_long2, P_long3, P_long4, P_long5, P_long6, P_long7, P_long8, P_long9, P_long10, P_long11, P_long12, P_long13, P_long14;


// Short D2S Conversion:

DEC2STCH D2S0(.CLK(CLK), .D(PD0), .LFSR(R0), .S(P0),.INIT(1'b0));
DEC2STCH D2S1(.CLK(CLK), .D(PD1), .LFSR(R1), .S(P1),.INIT(1'b0));
DEC2STCH D2S2(.CLK(CLK), .D(PD2), .LFSR(R2), .S(P2),.INIT(1'b0));
DEC2STCH D2S3(.CLK(CLK), .D(PD3), .LFSR(R3), .S(P3),.INIT(1'b0));
DEC2STCH D2S4(.CLK(CLK), .D(PD4), .LFSR(R4), .S(P4),.INIT(1'b0));
DEC2STCH D2S5(.CLK(CLK), .D(PD5), .LFSR(R5), .S(P5),.INIT(1'b0));
DEC2STCH D2S6(.CLK(CLK), .D(PD6), .LFSR(R6), .S(P6),.INIT(1'b0));
DEC2STCH D2S7(.CLK(CLK), .D(PD7), .LFSR(R7), .S(P7),.INIT(1'b0));
DEC2STCH D2S8(.CLK(CLK), .D(PD8), .LFSR(R8), .S(P8),.INIT(1'b0));
DEC2STCH D2S9(.CLK(CLK), .D(PD9), .LFSR(R9), .S(P9),.INIT(1'b0));
DEC2STCH D2S10(.CLK(CLK), .D(PD10), .LFSR(R10), .S(P10),.INIT(1'b0));
DEC2STCH D2S11(.CLK(CLK), .D(PD11), .LFSR(R11), .S(P11),.INIT(1'b0));
DEC2STCH D2S12(.CLK(CLK), .D(PD12), .LFSR(R12), .S(P12),.INIT(1'b0));
DEC2STCH D2S13(.CLK(CLK), .D(PD13), .LFSR(R13), .S(P13),.INIT(1'b0));
DEC2STCH D2S14(.CLK(CLK), .D(PD14), .LFSR(R14), .S(P14),.INIT(1'b0));
DEC2STCH D2S15(.CLK(CLK), .D(PD15), .LFSR(R15), .S(P15),.INIT(1'b0));
DEC2STCH D2S16(.CLK(CLK), .D(PD16), .LFSR(R16), .S(P16),.INIT(1'b0));
DEC2STCH D2S17(.CLK(CLK), .D(PD17), .LFSR(R17), .S(P17),.INIT(1'b0));
DEC2STCH D2S18(.CLK(CLK), .D(PD18), .LFSR(R18), .S(P18),.INIT(1'b0));
DEC2STCH D2S19(.CLK(CLK), .D(PD19), .LFSR(R19), .S(P19),.INIT(1'b0));
DEC2STCH D2S20(.CLK(CLK), .D(PD20), .LFSR(R20), .S(P20),.INIT(1'b0));
DEC2STCH D2S21(.CLK(CLK), .D(PD21), .LFSR(R21), .S(P21),.INIT(1'b0));
DEC2STCH D2S22(.CLK(CLK), .D(PD22), .LFSR(R22), .S(P22),.INIT(1'b0));
DEC2STCH D2S23(.CLK(CLK), .D(PD23), .LFSR(R23), .S(P23),.INIT(1'b0));
DEC2STCH D2S24(.CLK(CLK), .D(PD24), .LFSR(R24), .S(P24),.INIT(1'b0));
DEC2STCH D2S25(.CLK(CLK), .D(PD25), .LFSR(R25), .S(P25),.INIT(1'b0));
DEC2STCH D2S26(.CLK(CLK), .D(PD26), .LFSR(R26), .S(P26),.INIT(1'b0));
DEC2STCH D2S27(.CLK(CLK), .D(PD27), .LFSR(R27), .S(P27),.INIT(1'b0));
DEC2STCH D2S28(.CLK(CLK), .D(PD28), .LFSR(R28), .S(P28),.INIT(1'b0));
DEC2STCH D2S29(.CLK(CLK), .D(PD29), .LFSR(R29), .S(P29),.INIT(1'b0));
DEC2STCH D2S30(.CLK(CLK), .D(PD30), .LFSR(R30), .S(P30),.INIT(1'b0));
DEC2STCH D2S31(.CLK(CLK), .D(PD31), .LFSR(R31), .S(P31),.INIT(1'b0));
DEC2STCH D2S32(.CLK(CLK), .D(PD32), .LFSR(R32), .S(P32),.INIT(1'b0));
DEC2STCH D2S33(.CLK(CLK), .D(PD33), .LFSR(R33), .S(P33),.INIT(1'b0));
DEC2STCH D2S34(.CLK(CLK), .D(PD34), .LFSR(R34), .S(P34),.INIT(1'b0));
DEC2STCH D2S35(.CLK(CLK), .D(PD35), .LFSR(R35), .S(P35),.INIT(1'b0));
DEC2STCH D2S36(.CLK(CLK), .D(PD36), .LFSR(R36), .S(P36),.INIT(1'b0));
DEC2STCH D2S37(.CLK(CLK), .D(PD37), .LFSR(R37), .S(P37),.INIT(1'b0));
DEC2STCH D2S38(.CLK(CLK), .D(PD38), .LFSR(R38), .S(P38),.INIT(1'b0));
DEC2STCH D2S39(.CLK(CLK), .D(PD39), .LFSR(R39), .S(P39),.INIT(1'b0));
DEC2STCH D2S40(.CLK(CLK), .D(PD40), .LFSR(R40), .S(P40),.INIT(1'b0));
DEC2STCH D2S41(.CLK(CLK), .D(PD41), .LFSR(R41), .S(P41),.INIT(1'b0));
DEC2STCH D2S42(.CLK(CLK), .D(PD42), .LFSR(R42), .S(P42),.INIT(1'b0));
DEC2STCH D2S43(.CLK(CLK), .D(PD43), .LFSR(R43), .S(P43),.INIT(1'b0));
DEC2STCH D2S44(.CLK(CLK), .D(PD44), .LFSR(R44), .S(P44),.INIT(1'b0));
DEC2STCH D2S45(.CLK(CLK), .D(PD45), .LFSR(R45), .S(P45),.INIT(1'b0));
DEC2STCH D2S46(.CLK(CLK), .D(PD46), .LFSR(R46), .S(P46),.INIT(1'b0));
DEC2STCH D2S47(.CLK(CLK), .D(PD47), .LFSR(R47), .S(P47),.INIT(1'b0));
DEC2STCH D2S48(.CLK(CLK), .D(PD48), .LFSR(R48), .S(P48),.INIT(1'b0));
DEC2STCH D2S49(.CLK(CLK), .D(PD49), .LFSR(R49), .S(P49),.INIT(1'b0));
DEC2STCH D2S50(.CLK(CLK), .D(PD50), .LFSR(R50), .S(P50),.INIT(1'b0));
DEC2STCH D2S51(.CLK(CLK), .D(PD51), .LFSR(R51), .S(P51),.INIT(1'b0));
DEC2STCH D2S52(.CLK(CLK), .D(PD52), .LFSR(R52), .S(P52),.INIT(1'b0));
DEC2STCH D2S53(.CLK(CLK), .D(PD53), .LFSR(R53), .S(P53),.INIT(1'b0));
DEC2STCH D2S54(.CLK(CLK), .D(PD54), .LFSR(R54), .S(P54),.INIT(1'b0));
DEC2STCH D2S55(.CLK(CLK), .D(PD55), .LFSR(R55), .S(P55),.INIT(1'b0));
DEC2STCH D2S56(.CLK(CLK), .D(PD56), .LFSR(R56), .S(P56),.INIT(1'b0));
DEC2STCH D2S57(.CLK(CLK), .D(PD57), .LFSR(R57), .S(P57),.INIT(1'b0));
DEC2STCH D2S58(.CLK(CLK), .D(PD58), .LFSR(R58), .S(P58),.INIT(1'b0));
DEC2STCH D2S59(.CLK(CLK), .D(PD59), .LFSR(R59), .S(P59),.INIT(1'b0));
DEC2STCH D2S60(.CLK(CLK), .D(PD60), .LFSR(R60), .S(P60),.INIT(1'b0));
DEC2STCH D2S61(.CLK(CLK), .D(PD61), .LFSR(R61), .S(P61),.INIT(1'b0));
DEC2STCH D2S62(.CLK(CLK), .D(PD62), .LFSR(R62), .S(P62),.INIT(1'b0));
DEC2STCH D2S63(.CLK(CLK), .D(PD63), .LFSR(R63), .S(P63),.INIT(1'b0));
DEC2STCH D2S64(.CLK(CLK), .D(PD64), .LFSR(R64), .S(P64),.INIT(1'b0));
DEC2STCH D2S65(.CLK(CLK), .D(PD65), .LFSR(R65), .S(P65),.INIT(1'b0));
DEC2STCH D2S66(.CLK(CLK), .D(PD66), .LFSR(R66), .S(P66),.INIT(1'b0));
DEC2STCH D2S67(.CLK(CLK), .D(PD67), .LFSR(R67), .S(P67),.INIT(1'b0));
DEC2STCH D2S68(.CLK(CLK), .D(PD68), .LFSR(R68), .S(P68),.INIT(1'b0));
DEC2STCH D2S69(.CLK(CLK), .D(PD69), .LFSR(R69), .S(P69),.INIT(1'b0));
DEC2STCH D2S70(.CLK(CLK), .D(PD70), .LFSR(R70), .S(P70),.INIT(1'b0));
DEC2STCH D2S71(.CLK(CLK), .D(PD71), .LFSR(R71), .S(P71),.INIT(1'b0));
DEC2STCH D2S72(.CLK(CLK), .D(PD72), .LFSR(R72), .S(P72),.INIT(1'b0));
DEC2STCH D2S73(.CLK(CLK), .D(PD73), .LFSR(R73), .S(P73),.INIT(1'b0));
DEC2STCH D2S74(.CLK(CLK), .D(PD74), .LFSR(R74), .S(P74),.INIT(1'b0));
DEC2STCH D2S75(.CLK(CLK), .D(PD75), .LFSR(R75), .S(P75),.INIT(1'b0));
DEC2STCH D2S76(.CLK(CLK), .D(PD76), .LFSR(R76), .S(P76),.INIT(1'b0));
DEC2STCH D2S77(.CLK(CLK), .D(PD77), .LFSR(R77), .S(P77),.INIT(1'b0));
DEC2STCH D2S78(.CLK(CLK), .D(PD78), .LFSR(R78), .S(P78),.INIT(1'b0));
DEC2STCH D2S79(.CLK(CLK), .D(PD79), .LFSR(R79), .S(P79),.INIT(1'b0));
DEC2STCH D2S80(.CLK(CLK), .D(PD80), .LFSR(R80), .S(P80),.INIT(1'b0));
DEC2STCH D2S81(.CLK(CLK), .D(PD81), .LFSR(R81), .S(P81),.INIT(1'b0));
DEC2STCH D2S82(.CLK(CLK), .D(PD82), .LFSR(R82), .S(P82),.INIT(1'b0));
DEC2STCH D2S83(.CLK(CLK), .D(PD83), .LFSR(R83), .S(P83),.INIT(1'b0));
DEC2STCH D2S84(.CLK(CLK), .D(PD84), .LFSR(R84), .S(P84),.INIT(1'b0));
DEC2STCH D2S85(.CLK(CLK), .D(PD85), .LFSR(R85), .S(P85),.INIT(1'b0));
DEC2STCH D2S86(.CLK(CLK), .D(PD86), .LFSR(R86), .S(P86),.INIT(1'b0));
DEC2STCH D2S87(.CLK(CLK), .D(PD87), .LFSR(R87), .S(P87),.INIT(1'b0));
DEC2STCH D2S88(.CLK(CLK), .D(PD88), .LFSR(R88), .S(P88),.INIT(1'b0));
DEC2STCH D2S89(.CLK(CLK), .D(PD89), .LFSR(R89), .S(P89),.INIT(1'b0));
DEC2STCH D2S90(.CLK(CLK), .D(PD90), .LFSR(R90), .S(P90),.INIT(1'b0));
DEC2STCH D2S91(.CLK(CLK), .D(PD91), .LFSR(R91), .S(P91),.INIT(1'b0));
DEC2STCH D2S92(.CLK(CLK), .D(PD92), .LFSR(R92), .S(P92),.INIT(1'b0));
DEC2STCH D2S93(.CLK(CLK), .D(PD93), .LFSR(R93), .S(P93),.INIT(1'b0));
DEC2STCH D2S94(.CLK(CLK), .D(PD94), .LFSR(R94), .S(P94),.INIT(1'b0));
DEC2STCH D2S95(.CLK(CLK), .D(PD95), .LFSR(R95), .S(P95),.INIT(1'b0));
DEC2STCH D2S96(.CLK(CLK), .D(PD96), .LFSR(R96), .S(P96),.INIT(1'b0));
DEC2STCH D2S97(.CLK(CLK), .D(PD97), .LFSR(R97), .S(P97),.INIT(1'b0));
DEC2STCH D2S98(.CLK(CLK), .D(PD98), .LFSR(R98), .S(P98),.INIT(1'b0));
DEC2STCH D2S99(.CLK(CLK), .D(PD99), .LFSR(R99), .S(P99),.INIT(1'b0));
DEC2STCH D2S100(.CLK(CLK), .D(PD100), .LFSR(R100), .S(P100),.INIT(1'b0));
DEC2STCH D2S101(.CLK(CLK), .D(PD101), .LFSR(R101), .S(P101),.INIT(1'b0));
DEC2STCH D2S102(.CLK(CLK), .D(PD102), .LFSR(R102), .S(P102),.INIT(1'b0));
DEC2STCH D2S103(.CLK(CLK), .D(PD103), .LFSR(R103), .S(P103),.INIT(1'b0));
DEC2STCH D2S104(.CLK(CLK), .D(PD104), .LFSR(R104), .S(P104),.INIT(1'b0));
DEC2STCH D2S105(.CLK(CLK), .D(PD105), .LFSR(R105), .S(P105),.INIT(1'b0));
DEC2STCH D2S106(.CLK(CLK), .D(PD106), .LFSR(R106), .S(P106),.INIT(1'b0));
DEC2STCH D2S107(.CLK(CLK), .D(PD107), .LFSR(R107), .S(P107),.INIT(1'b0));
DEC2STCH D2S108(.CLK(CLK), .D(PD108), .LFSR(R108), .S(P108),.INIT(1'b0));
DEC2STCH D2S109(.CLK(CLK), .D(PD109), .LFSR(R109), .S(P109),.INIT(1'b0));
DEC2STCH D2S110(.CLK(CLK), .D(PD110), .LFSR(R110), .S(P110),.INIT(1'b0));
DEC2STCH D2S111(.CLK(CLK), .D(PD111), .LFSR(R111), .S(P111),.INIT(1'b0));
DEC2STCH D2S112(.CLK(CLK), .D(PD112), .LFSR(R112), .S(P112),.INIT(1'b0));
DEC2STCH D2S113(.CLK(CLK), .D(PD113), .LFSR(R113), .S(P113),.INIT(1'b0));
DEC2STCH D2S114(.CLK(CLK), .D(PD114), .LFSR(R114), .S(P114),.INIT(1'b0));
DEC2STCH D2S115(.CLK(CLK), .D(PD115), .LFSR(R115), .S(P115),.INIT(1'b0));
DEC2STCH D2S116(.CLK(CLK), .D(PD116), .LFSR(R116), .S(P116),.INIT(1'b0));
DEC2STCH D2S117(.CLK(CLK), .D(PD117), .LFSR(R117), .S(P117),.INIT(1'b0));
DEC2STCH D2S118(.CLK(CLK), .D(PD118), .LFSR(R118), .S(P118),.INIT(1'b0));
DEC2STCH D2S119(.CLK(CLK), .D(PD119), .LFSR(R119), .S(P119),.INIT(1'b0));
DEC2STCH D2S120(.CLK(CLK), .D(PD120), .LFSR(R120), .S(P120),.INIT(1'b0));
DEC2STCH D2S121(.CLK(CLK), .D(PD121), .LFSR(R121), .S(P121),.INIT(1'b0));
DEC2STCH D2S122(.CLK(CLK), .D(PD122), .LFSR(R122), .S(P122),.INIT(1'b0));
DEC2STCH D2S123(.CLK(CLK), .D(PD123), .LFSR(R123), .S(P123),.INIT(1'b0));
DEC2STCH D2S124(.CLK(CLK), .D(PD124), .LFSR(R124), .S(P124),.INIT(1'b0));
DEC2STCH D2S125(.CLK(CLK), .D(PD125), .LFSR(R125), .S(P125),.INIT(1'b0));
DEC2STCH D2S126(.CLK(CLK), .D(PD126), .LFSR(R126), .S(P126),.INIT(1'b0));
DEC2STCH D2S127(.CLK(CLK), .D(PD127), .LFSR(R127), .S(P127),.INIT(1'b0));
DEC2STCH D2S128(.CLK(CLK), .D(PD128), .LFSR(R128), .S(P128),.INIT(1'b0));
DEC2STCH D2S129(.CLK(CLK), .D(PD129), .LFSR(R129), .S(P129),.INIT(1'b0));
DEC2STCH D2S130(.CLK(CLK), .D(PD130), .LFSR(R130), .S(P130),.INIT(1'b0));
DEC2STCH D2S131(.CLK(CLK), .D(PD131), .LFSR(R131), .S(P131),.INIT(1'b0));
DEC2STCH D2S132(.CLK(CLK), .D(PD132), .LFSR(R132), .S(P132),.INIT(1'b0));
DEC2STCH D2S133(.CLK(CLK), .D(PD133), .LFSR(R133), .S(P133),.INIT(1'b0));
DEC2STCH D2S134(.CLK(CLK), .D(PD134), .LFSR(R134), .S(P134),.INIT(1'b0));
DEC2STCH D2S135(.CLK(CLK), .D(PD135), .LFSR(R135), .S(P135),.INIT(1'b0));
DEC2STCH D2S136(.CLK(CLK), .D(PD136), .LFSR(R136), .S(P136),.INIT(1'b0));
DEC2STCH D2S137(.CLK(CLK), .D(PD137), .LFSR(R137), .S(P137),.INIT(1'b0));
DEC2STCH D2S138(.CLK(CLK), .D(PD138), .LFSR(R138), .S(P138),.INIT(1'b0));
DEC2STCH D2S139(.CLK(CLK), .D(PD139), .LFSR(R139), .S(P139),.INIT(1'b0));
DEC2STCH D2S140(.CLK(CLK), .D(PD140), .LFSR(R140), .S(P140),.INIT(1'b0));
DEC2STCH D2S141(.CLK(CLK), .D(PD141), .LFSR(R141), .S(P141),.INIT(1'b0));
DEC2STCH D2S142(.CLK(CLK), .D(PD142), .LFSR(R142), .S(P142),.INIT(1'b0));
DEC2STCH D2S143(.CLK(CLK), .D(PD143), .LFSR(R143), .S(P143),.INIT(1'b0));
DEC2STCH D2S144(.CLK(CLK), .D(PD144), .LFSR(R144), .S(P144),.INIT(1'b0));
DEC2STCH D2S145(.CLK(CLK), .D(PD145), .LFSR(R145), .S(P145),.INIT(1'b0));
DEC2STCH D2S146(.CLK(CLK), .D(PD146), .LFSR(R146), .S(P146),.INIT(1'b0));
DEC2STCH D2S147(.CLK(CLK), .D(PD147), .LFSR(R147), .S(P147),.INIT(1'b0));
DEC2STCH D2S148(.CLK(CLK), .D(PD148), .LFSR(R148), .S(P148),.INIT(1'b0));
DEC2STCH D2S149(.CLK(CLK), .D(PD149), .LFSR(R149), .S(P149),.INIT(1'b0));
DEC2STCH D2S150(.CLK(CLK), .D(PD150), .LFSR(R150), .S(P150),.INIT(1'b0));
DEC2STCH D2S151(.CLK(CLK), .D(PD151), .LFSR(R151), .S(P151),.INIT(1'b0));
DEC2STCH D2S152(.CLK(CLK), .D(PD152), .LFSR(R152), .S(P152),.INIT(1'b0));
DEC2STCH D2S153(.CLK(CLK), .D(PD153), .LFSR(R153), .S(P153),.INIT(1'b0));
DEC2STCH D2S154(.CLK(CLK), .D(PD154), .LFSR(R154), .S(P154),.INIT(1'b0));
DEC2STCH D2S155(.CLK(CLK), .D(PD155), .LFSR(R155), .S(P155),.INIT(1'b0));
DEC2STCH D2S156(.CLK(CLK), .D(PD156), .LFSR(R156), .S(P156),.INIT(1'b0));
DEC2STCH D2S157(.CLK(CLK), .D(PD157), .LFSR(R157), .S(P157),.INIT(1'b0));
DEC2STCH D2S158(.CLK(CLK), .D(PD158), .LFSR(R158), .S(P158),.INIT(1'b0));
DEC2STCH D2S159(.CLK(CLK), .D(PD159), .LFSR(R159), .S(P159),.INIT(1'b0));
DEC2STCH D2S160(.CLK(CLK), .D(PD160), .LFSR(R160), .S(P160),.INIT(1'b0));
DEC2STCH D2S161(.CLK(CLK), .D(PD161), .LFSR(R161), .S(P161),.INIT(1'b0));
DEC2STCH D2S162(.CLK(CLK), .D(PD162), .LFSR(R162), .S(P162),.INIT(1'b0));
DEC2STCH D2S163(.CLK(CLK), .D(PD163), .LFSR(R163), .S(P163),.INIT(1'b0));
DEC2STCH D2S164(.CLK(CLK), .D(PD164), .LFSR(R164), .S(P164),.INIT(1'b0));
DEC2STCH D2S165(.CLK(CLK), .D(PD165), .LFSR(R165), .S(P165),.INIT(1'b0));
DEC2STCH D2S166(.CLK(CLK), .D(PD166), .LFSR(R166), .S(P166),.INIT(1'b0));
DEC2STCH D2S167(.CLK(CLK), .D(PD167), .LFSR(R167), .S(P167),.INIT(1'b0));
DEC2STCH D2S168(.CLK(CLK), .D(PD168), .LFSR(R168), .S(P168),.INIT(1'b0));
DEC2STCH D2S169(.CLK(CLK), .D(PD169), .LFSR(R169), .S(P169),.INIT(1'b0));
DEC2STCH D2S170(.CLK(CLK), .D(PD170), .LFSR(R170), .S(P170),.INIT(1'b0));
DEC2STCH D2S171(.CLK(CLK), .D(PD171), .LFSR(R171), .S(P171),.INIT(1'b0));
DEC2STCH D2S172(.CLK(CLK), .D(PD172), .LFSR(R172), .S(P172),.INIT(1'b0));
DEC2STCH D2S173(.CLK(CLK), .D(PD173), .LFSR(R173), .S(P173),.INIT(1'b0));
DEC2STCH D2S174(.CLK(CLK), .D(PD174), .LFSR(R174), .S(P174),.INIT(1'b0));
DEC2STCH D2S175(.CLK(CLK), .D(PD175), .LFSR(R175), .S(P175),.INIT(1'b0));
DEC2STCH D2S176(.CLK(CLK), .D(PD176), .LFSR(R176), .S(P176),.INIT(1'b0));
DEC2STCH D2S177(.CLK(CLK), .D(PD177), .LFSR(R177), .S(P177),.INIT(1'b0));
DEC2STCH D2S178(.CLK(CLK), .D(PD178), .LFSR(R178), .S(P178),.INIT(1'b0));
DEC2STCH D2S179(.CLK(CLK), .D(PD179), .LFSR(R179), .S(P179),.INIT(1'b0));
DEC2STCH D2S180(.CLK(CLK), .D(PD180), .LFSR(R180), .S(P180),.INIT(1'b0));
DEC2STCH D2S181(.CLK(CLK), .D(PD181), .LFSR(R181), .S(P181),.INIT(1'b0));
DEC2STCH D2S182(.CLK(CLK), .D(PD182), .LFSR(R182), .S(P182),.INIT(1'b0));
DEC2STCH D2S183(.CLK(CLK), .D(PD183), .LFSR(R183), .S(P183),.INIT(1'b0));
DEC2STCH D2S184(.CLK(CLK), .D(PD184), .LFSR(R184), .S(P184),.INIT(1'b0));
DEC2STCH D2S185(.CLK(CLK), .D(PD185), .LFSR(R185), .S(P185),.INIT(1'b0));
DEC2STCH D2S186(.CLK(CLK), .D(PD186), .LFSR(R186), .S(P186),.INIT(1'b0));
DEC2STCH D2S187(.CLK(CLK), .D(PD187), .LFSR(R187), .S(P187),.INIT(1'b0));
DEC2STCH D2S188(.CLK(CLK), .D(PD188), .LFSR(R188), .S(P188),.INIT(1'b0));
DEC2STCH D2S189(.CLK(CLK), .D(PD189), .LFSR(R189), .S(P189),.INIT(1'b0));
DEC2STCH D2S190(.CLK(CLK), .D(PD190), .LFSR(R190), .S(P190),.INIT(1'b0));
DEC2STCH D2S191(.CLK(CLK), .D(PD191), .LFSR(R191), .S(P191),.INIT(1'b0));
DEC2STCH D2S192(.CLK(CLK), .D(PD192), .LFSR(R192), .S(P192),.INIT(1'b0));
DEC2STCH D2S193(.CLK(CLK), .D(PD193), .LFSR(R193), .S(P193),.INIT(1'b0));
DEC2STCH D2S194(.CLK(CLK), .D(PD194), .LFSR(R194), .S(P194),.INIT(1'b0));
DEC2STCH D2S195(.CLK(CLK), .D(PD195), .LFSR(R195), .S(P195),.INIT(1'b0));
DEC2STCH D2S196(.CLK(CLK), .D(PD196), .LFSR(R196), .S(P196),.INIT(1'b0));
DEC2STCH D2S197(.CLK(CLK), .D(PD197), .LFSR(R197), .S(P197),.INIT(1'b0));
DEC2STCH D2S198(.CLK(CLK), .D(PD198), .LFSR(R198), .S(P198),.INIT(1'b0));
DEC2STCH D2S199(.CLK(CLK), .D(PD199), .LFSR(R199), .S(P199),.INIT(1'b0));
DEC2STCH D2S200(.CLK(CLK), .D(PD200), .LFSR(R200), .S(P200),.INIT(1'b0));
DEC2STCH D2S201(.CLK(CLK), .D(PD201), .LFSR(R201), .S(P201),.INIT(1'b0));
DEC2STCH D2S202(.CLK(CLK), .D(PD202), .LFSR(R202), .S(P202),.INIT(1'b0));
DEC2STCH D2S203(.CLK(CLK), .D(PD203), .LFSR(R203), .S(P203),.INIT(1'b0));
DEC2STCH D2S204(.CLK(CLK), .D(PD204), .LFSR(R204), .S(P204),.INIT(1'b0));
DEC2STCH D2S205(.CLK(CLK), .D(PD205), .LFSR(R205), .S(P205),.INIT(1'b0));
DEC2STCH D2S206(.CLK(CLK), .D(PD206), .LFSR(R206), .S(P206),.INIT(1'b0));
DEC2STCH D2S207(.CLK(CLK), .D(PD207), .LFSR(R207), .S(P207),.INIT(1'b0));
DEC2STCH D2S208(.CLK(CLK), .D(PD208), .LFSR(R208), .S(P208),.INIT(1'b0));
DEC2STCH D2S209(.CLK(CLK), .D(PD209), .LFSR(R209), .S(P209),.INIT(1'b0));
DEC2STCH D2S210(.CLK(CLK), .D(PD210), .LFSR(R210), .S(P210),.INIT(1'b0));
DEC2STCH D2S211(.CLK(CLK), .D(PD211), .LFSR(R211), .S(P211),.INIT(1'b0));
DEC2STCH D2S212(.CLK(CLK), .D(PD212), .LFSR(R212), .S(P212),.INIT(1'b0));
DEC2STCH D2S213(.CLK(CLK), .D(PD213), .LFSR(R213), .S(P213),.INIT(1'b0));
DEC2STCH D2S214(.CLK(CLK), .D(PD214), .LFSR(R214), .S(P214),.INIT(1'b0));
DEC2STCH D2S215(.CLK(CLK), .D(PD215), .LFSR(R215), .S(P215),.INIT(1'b0));
DEC2STCH D2S216(.CLK(CLK), .D(PD216), .LFSR(R216), .S(P216),.INIT(1'b0));
DEC2STCH D2S217(.CLK(CLK), .D(PD217), .LFSR(R217), .S(P217),.INIT(1'b0));
DEC2STCH D2S218(.CLK(CLK), .D(PD218), .LFSR(R218), .S(P218),.INIT(1'b0));
DEC2STCH D2S219(.CLK(CLK), .D(PD219), .LFSR(R219), .S(P219),.INIT(1'b0));
DEC2STCH D2S220(.CLK(CLK), .D(PD220), .LFSR(R220), .S(P220),.INIT(1'b0));
DEC2STCH D2S221(.CLK(CLK), .D(PD221), .LFSR(R221), .S(P221),.INIT(1'b0));
DEC2STCH D2S222(.CLK(CLK), .D(PD222), .LFSR(R222), .S(P222),.INIT(1'b0));
DEC2STCH D2S223(.CLK(CLK), .D(PD223), .LFSR(R223), .S(P223),.INIT(1'b0));
DEC2STCH D2S224(.CLK(CLK), .D(PD224), .LFSR(R224), .S(P224),.INIT(1'b0));
DEC2STCH D2S225(.CLK(CLK), .D(PD225), .LFSR(R225), .S(P225),.INIT(1'b0));
DEC2STCH D2S226(.CLK(CLK), .D(PD226), .LFSR(R226), .S(P226),.INIT(1'b0));
DEC2STCH D2S227(.CLK(CLK), .D(PD227), .LFSR(R227), .S(P227),.INIT(1'b0));
DEC2STCH D2S228(.CLK(CLK), .D(PD228), .LFSR(R228), .S(P228),.INIT(1'b0));
DEC2STCH D2S229(.CLK(CLK), .D(PD229), .LFSR(R229), .S(P229),.INIT(1'b0));
DEC2STCH D2S230(.CLK(CLK), .D(PD230), .LFSR(R230), .S(P230),.INIT(1'b0));
DEC2STCH D2S231(.CLK(CLK), .D(PD231), .LFSR(R231), .S(P231),.INIT(1'b0));
DEC2STCH D2S232(.CLK(CLK), .D(PD232), .LFSR(R232), .S(P232),.INIT(1'b0));
DEC2STCH D2S233(.CLK(CLK), .D(PD233), .LFSR(R233), .S(P233),.INIT(1'b0));
DEC2STCH D2S234(.CLK(CLK), .D(PD234), .LFSR(R234), .S(P234),.INIT(1'b0));
DEC2STCH D2S235(.CLK(CLK), .D(PD235), .LFSR(R235), .S(P235),.INIT(1'b0));
DEC2STCH D2S236(.CLK(CLK), .D(PD236), .LFSR(R236), .S(P236),.INIT(1'b0));
DEC2STCH D2S237(.CLK(CLK), .D(PD237), .LFSR(R237), .S(P237),.INIT(1'b0));
DEC2STCH D2S238(.CLK(CLK), .D(PD238), .LFSR(R238), .S(P238),.INIT(1'b0));
DEC2STCH D2S239(.CLK(CLK), .D(PD239), .LFSR(R239), .S(P239),.INIT(1'b0));
DEC2STCH D2S240(.CLK(CLK), .D(PD240), .LFSR(R240), .S(P240),.INIT(1'b0));
DEC2STCH D2S241(.CLK(CLK), .D(PD241), .LFSR(R241), .S(P241),.INIT(1'b0));
DEC2STCH D2S242(.CLK(CLK), .D(PD242), .LFSR(R242), .S(P242),.INIT(1'b0));
DEC2STCH D2S243(.CLK(CLK), .D(PD243), .LFSR(R243), .S(P243),.INIT(1'b0));
DEC2STCH D2S244(.CLK(CLK), .D(PD244), .LFSR(R244), .S(P244),.INIT(1'b0));
DEC2STCH D2S245(.CLK(CLK), .D(PD245), .LFSR(R245), .S(P245),.INIT(1'b0));
DEC2STCH D2S246(.CLK(CLK), .D(PD246), .LFSR(R246), .S(P246),.INIT(1'b0));
DEC2STCH D2S247(.CLK(CLK), .D(PD247), .LFSR(R247), .S(P247),.INIT(1'b0));
DEC2STCH D2S248(.CLK(CLK), .D(PD248), .LFSR(R248), .S(P248),.INIT(1'b0));
DEC2STCH D2S249(.CLK(CLK), .D(PD249), .LFSR(R249), .S(P249),.INIT(1'b0));
DEC2STCH D2S250(.CLK(CLK), .D(PD250), .LFSR(R250), .S(P250),.INIT(1'b0));
DEC2STCH D2S251(.CLK(CLK), .D(PD251), .LFSR(R251), .S(P251),.INIT(1'b0));
DEC2STCH D2S252(.CLK(CLK), .D(PD252), .LFSR(R252), .S(P252),.INIT(1'b0));
DEC2STCH D2S253(.CLK(CLK), .D(PD253), .LFSR(R253), .S(P253),.INIT(1'b0));
DEC2STCH D2S254(.CLK(CLK), .D(PD254), .LFSR(R254), .S(P254),.INIT(1'b0));
DEC2STCH D2S255(.CLK(CLK), .D(PD255), .LFSR(R255), .S(P255),.INIT(1'b0));
DEC2STCH D2S256(.CLK(CLK), .D(PD256), .LFSR(R256), .S(P256),.INIT(1'b0));
DEC2STCH D2S257(.CLK(CLK), .D(PD257), .LFSR(R257), .S(P257),.INIT(1'b0));
DEC2STCH D2S258(.CLK(CLK), .D(PD258), .LFSR(R258), .S(P258),.INIT(1'b0));
DEC2STCH D2S259(.CLK(CLK), .D(PD259), .LFSR(R259), .S(P259),.INIT(1'b0));
DEC2STCH D2S260(.CLK(CLK), .D(PD260), .LFSR(R260), .S(P260),.INIT(1'b0));
DEC2STCH D2S261(.CLK(CLK), .D(PD261), .LFSR(R261), .S(P261),.INIT(1'b0));
DEC2STCH D2S262(.CLK(CLK), .D(PD262), .LFSR(R262), .S(P262),.INIT(1'b0));
DEC2STCH D2S263(.CLK(CLK), .D(PD263), .LFSR(R263), .S(P263),.INIT(1'b0));
DEC2STCH D2S264(.CLK(CLK), .D(PD264), .LFSR(R264), .S(P264),.INIT(1'b0));
DEC2STCH D2S265(.CLK(CLK), .D(PD265), .LFSR(R265), .S(P265),.INIT(1'b0));
DEC2STCH D2S266(.CLK(CLK), .D(PD266), .LFSR(R266), .S(P266),.INIT(1'b0));
DEC2STCH D2S267(.CLK(CLK), .D(PD267), .LFSR(R267), .S(P267),.INIT(1'b0));
DEC2STCH D2S268(.CLK(CLK), .D(PD268), .LFSR(R268), .S(P268),.INIT(1'b0));
DEC2STCH D2S269(.CLK(CLK), .D(PD269), .LFSR(R269), .S(P269),.INIT(1'b0));
DEC2STCH D2S270(.CLK(CLK), .D(PD270), .LFSR(R270), .S(P270),.INIT(1'b0));
DEC2STCH D2S271(.CLK(CLK), .D(PD271), .LFSR(R271), .S(P271),.INIT(1'b0));
DEC2STCH D2S272(.CLK(CLK), .D(PD272), .LFSR(R272), .S(P272),.INIT(1'b0));
DEC2STCH D2S273(.CLK(CLK), .D(PD273), .LFSR(R273), .S(P273),.INIT(1'b0));
DEC2STCH D2S274(.CLK(CLK), .D(PD274), .LFSR(R274), .S(P274),.INIT(1'b0));
DEC2STCH D2S275(.CLK(CLK), .D(PD275), .LFSR(R275), .S(P275),.INIT(1'b0));
DEC2STCH D2S276(.CLK(CLK), .D(PD276), .LFSR(R276), .S(P276),.INIT(1'b0));
DEC2STCH D2S277(.CLK(CLK), .D(PD277), .LFSR(R277), .S(P277),.INIT(1'b0));
DEC2STCH D2S278(.CLK(CLK), .D(PD278), .LFSR(R278), .S(P278),.INIT(1'b0));
DEC2STCH D2S279(.CLK(CLK), .D(PD279), .LFSR(R279), .S(P279),.INIT(1'b0));
DEC2STCH D2S280(.CLK(CLK), .D(PD280), .LFSR(R280), .S(P280),.INIT(1'b0));
DEC2STCH D2S281(.CLK(CLK), .D(PD281), .LFSR(R281), .S(P281),.INIT(1'b0));
DEC2STCH D2S282(.CLK(CLK), .D(PD282), .LFSR(R282), .S(P282),.INIT(1'b0));
DEC2STCH D2S283(.CLK(CLK), .D(PD283), .LFSR(R283), .S(P283),.INIT(1'b0));
DEC2STCH D2S284(.CLK(CLK), .D(PD284), .LFSR(R284), .S(P284),.INIT(1'b0));
DEC2STCH D2S285(.CLK(CLK), .D(PD285), .LFSR(R285), .S(P285),.INIT(1'b0));
DEC2STCH D2S286(.CLK(CLK), .D(PD286), .LFSR(R286), .S(P286),.INIT(1'b0));
DEC2STCH D2S287(.CLK(CLK), .D(PD287), .LFSR(R287), .S(P287),.INIT(1'b0));
DEC2STCH D2S288(.CLK(CLK), .D(PD288), .LFSR(R288), .S(P288),.INIT(1'b0));
DEC2STCH D2S289(.CLK(CLK), .D(PD289), .LFSR(R289), .S(P289),.INIT(1'b0));
DEC2STCH D2S290(.CLK(CLK), .D(PD290), .LFSR(R290), .S(P290),.INIT(1'b0));
DEC2STCH D2S291(.CLK(CLK), .D(PD291), .LFSR(R291), .S(P291),.INIT(1'b0));
DEC2STCH D2S292(.CLK(CLK), .D(PD292), .LFSR(R292), .S(P292),.INIT(1'b0));
DEC2STCH D2S293(.CLK(CLK), .D(PD293), .LFSR(R293), .S(P293),.INIT(1'b0));
DEC2STCH D2S294(.CLK(CLK), .D(PD294), .LFSR(R294), .S(P294),.INIT(1'b0));
DEC2STCH D2S295(.CLK(CLK), .D(PD295), .LFSR(R295), .S(P295),.INIT(1'b0));
DEC2STCH D2S296(.CLK(CLK), .D(PD296), .LFSR(R296), .S(P296),.INIT(1'b0));
DEC2STCH D2S297(.CLK(CLK), .D(PD297), .LFSR(R297), .S(P297),.INIT(1'b0));
DEC2STCH D2S298(.CLK(CLK), .D(PD298), .LFSR(R298), .S(P298),.INIT(1'b0));
DEC2STCH D2S299(.CLK(CLK), .D(PD299), .LFSR(R299), .S(P299),.INIT(1'b0));
DEC2STCH D2S300(.CLK(CLK), .D(PD300), .LFSR(R300), .S(P300),.INIT(1'b0));
DEC2STCH D2S301(.CLK(CLK), .D(PD301), .LFSR(R301), .S(P301),.INIT(1'b0));
DEC2STCH D2S302(.CLK(CLK), .D(PD302), .LFSR(R302), .S(P302),.INIT(1'b0));
DEC2STCH D2S303(.CLK(CLK), .D(PD303), .LFSR(R303), .S(P303),.INIT(1'b0));
DEC2STCH D2S304(.CLK(CLK), .D(PD304), .LFSR(R304), .S(P304),.INIT(1'b0));
DEC2STCH D2S305(.CLK(CLK), .D(PD305), .LFSR(R305), .S(P305),.INIT(1'b0));
DEC2STCH D2S306(.CLK(CLK), .D(PD306), .LFSR(R306), .S(P306),.INIT(1'b0));
DEC2STCH D2S307(.CLK(CLK), .D(PD307), .LFSR(R307), .S(P307),.INIT(1'b0));
DEC2STCH D2S308(.CLK(CLK), .D(PD308), .LFSR(R308), .S(P308),.INIT(1'b0));
DEC2STCH D2S309(.CLK(CLK), .D(PD309), .LFSR(R309), .S(P309),.INIT(1'b0));
DEC2STCH D2S310(.CLK(CLK), .D(PD310), .LFSR(R310), .S(P310),.INIT(1'b0));
DEC2STCH D2S311(.CLK(CLK), .D(PD311), .LFSR(R311), .S(P311),.INIT(1'b0));
DEC2STCH D2S312(.CLK(CLK), .D(PD312), .LFSR(R312), .S(P312),.INIT(1'b0));
DEC2STCH D2S313(.CLK(CLK), .D(PD313), .LFSR(R313), .S(P313),.INIT(1'b0));
DEC2STCH D2S314(.CLK(CLK), .D(PD314), .LFSR(R314), .S(P314),.INIT(1'b0));
DEC2STCH D2S315(.CLK(CLK), .D(PD315), .LFSR(R315), .S(P315),.INIT(1'b0));
DEC2STCH D2S316(.CLK(CLK), .D(PD316), .LFSR(R316), .S(P316),.INIT(1'b0));
DEC2STCH D2S317(.CLK(CLK), .D(PD317), .LFSR(R317), .S(P317),.INIT(1'b0));
DEC2STCH D2S318(.CLK(CLK), .D(PD318), .LFSR(R318), .S(P318),.INIT(1'b0));
DEC2STCH D2S319(.CLK(CLK), .D(PD319), .LFSR(R319), .S(P319),.INIT(1'b0));
DEC2STCH D2S320(.CLK(CLK), .D(PD320), .LFSR(R320), .S(P320),.INIT(1'b0));
DEC2STCH D2S321(.CLK(CLK), .D(PD321), .LFSR(R321), .S(P321),.INIT(1'b0));
DEC2STCH D2S322(.CLK(CLK), .D(PD322), .LFSR(R322), .S(P322),.INIT(1'b0));
DEC2STCH D2S323(.CLK(CLK), .D(PD323), .LFSR(R323), .S(P323),.INIT(1'b0));
DEC2STCH D2S324(.CLK(CLK), .D(PD324), .LFSR(R324), .S(P324),.INIT(1'b0));
DEC2STCH D2S325(.CLK(CLK), .D(PD325), .LFSR(R325), .S(P325),.INIT(1'b0));
DEC2STCH D2S326(.CLK(CLK), .D(PD326), .LFSR(R326), .S(P326),.INIT(1'b0));
DEC2STCH D2S327(.CLK(CLK), .D(PD327), .LFSR(R327), .S(P327),.INIT(1'b0));
DEC2STCH D2S328(.CLK(CLK), .D(PD328), .LFSR(R328), .S(P328),.INIT(1'b0));
DEC2STCH D2S329(.CLK(CLK), .D(PD329), .LFSR(R329), .S(P329),.INIT(1'b0));
DEC2STCH D2S330(.CLK(CLK), .D(PD330), .LFSR(R330), .S(P330),.INIT(1'b0));
DEC2STCH D2S331(.CLK(CLK), .D(PD331), .LFSR(R331), .S(P331),.INIT(1'b0));
DEC2STCH D2S332(.CLK(CLK), .D(PD332), .LFSR(R332), .S(P332),.INIT(1'b0));
DEC2STCH D2S333(.CLK(CLK), .D(PD333), .LFSR(R333), .S(P333),.INIT(1'b0));
DEC2STCH D2S334(.CLK(CLK), .D(PD334), .LFSR(R334), .S(P334),.INIT(1'b0));
DEC2STCH D2S335(.CLK(CLK), .D(PD335), .LFSR(R335), .S(P335),.INIT(1'b0));
DEC2STCH D2S336(.CLK(CLK), .D(PD336), .LFSR(R336), .S(P336),.INIT(1'b0));
DEC2STCH D2S337(.CLK(CLK), .D(PD337), .LFSR(R337), .S(P337),.INIT(1'b0));
DEC2STCH D2S338(.CLK(CLK), .D(PD338), .LFSR(R338), .S(P338),.INIT(1'b0));
DEC2STCH D2S339(.CLK(CLK), .D(PD339), .LFSR(R339), .S(P339),.INIT(1'b0));
DEC2STCH D2S340(.CLK(CLK), .D(PD340), .LFSR(R340), .S(P340),.INIT(1'b0));
DEC2STCH D2S341(.CLK(CLK), .D(PD341), .LFSR(R341), .S(P341),.INIT(1'b0));
DEC2STCH D2S342(.CLK(CLK), .D(PD342), .LFSR(R342), .S(P342),.INIT(1'b0));
DEC2STCH D2S343(.CLK(CLK), .D(PD343), .LFSR(R343), .S(P343),.INIT(1'b0));
DEC2STCH D2S344(.CLK(CLK), .D(PD344), .LFSR(R344), .S(P344),.INIT(1'b0));
DEC2STCH D2S345(.CLK(CLK), .D(PD345), .LFSR(R345), .S(P345),.INIT(1'b0));
DEC2STCH D2S346(.CLK(CLK), .D(PD346), .LFSR(R346), .S(P346),.INIT(1'b0));
DEC2STCH D2S347(.CLK(CLK), .D(PD347), .LFSR(R347), .S(P347),.INIT(1'b0));
DEC2STCH D2S348(.CLK(CLK), .D(PD348), .LFSR(R348), .S(P348),.INIT(1'b0));
DEC2STCH D2S349(.CLK(CLK), .D(PD349), .LFSR(R349), .S(P349),.INIT(1'b0));
DEC2STCH D2S350(.CLK(CLK), .D(PD350), .LFSR(R350), .S(P350),.INIT(1'b0));
DEC2STCH D2S351(.CLK(CLK), .D(PD351), .LFSR(R351), .S(P351),.INIT(1'b0));
DEC2STCH D2S352(.CLK(CLK), .D(PD352), .LFSR(R352), .S(P352),.INIT(1'b0));
DEC2STCH D2S353(.CLK(CLK), .D(PD353), .LFSR(R353), .S(P353),.INIT(1'b0));
DEC2STCH D2S354(.CLK(CLK), .D(PD354), .LFSR(R354), .S(P354),.INIT(1'b0));
DEC2STCH D2S355(.CLK(CLK), .D(PD355), .LFSR(R355), .S(P355),.INIT(1'b0));
DEC2STCH D2S356(.CLK(CLK), .D(PD356), .LFSR(R356), .S(P356),.INIT(1'b0));
DEC2STCH D2S357(.CLK(CLK), .D(PD357), .LFSR(R357), .S(P357),.INIT(1'b0));
DEC2STCH D2S358(.CLK(CLK), .D(PD358), .LFSR(R358), .S(P358),.INIT(1'b0));
DEC2STCH D2S359(.CLK(CLK), .D(PD359), .LFSR(R359), .S(P359),.INIT(1'b0));
DEC2STCH D2S360(.CLK(CLK), .D(PD360), .LFSR(R360), .S(P360),.INIT(1'b0));
DEC2STCH D2S361(.CLK(CLK), .D(PD361), .LFSR(R361), .S(P361),.INIT(1'b0));
DEC2STCH D2S362(.CLK(CLK), .D(PD362), .LFSR(R362), .S(P362),.INIT(1'b0));
DEC2STCH D2S363(.CLK(CLK), .D(PD363), .LFSR(R363), .S(P363),.INIT(1'b0));
DEC2STCH D2S364(.CLK(CLK), .D(PD364), .LFSR(R364), .S(P364),.INIT(1'b0));
DEC2STCH D2S365(.CLK(CLK), .D(PD365), .LFSR(R365), .S(P365),.INIT(1'b0));
DEC2STCH D2S366(.CLK(CLK), .D(PD366), .LFSR(R366), .S(P366),.INIT(1'b0));
DEC2STCH D2S367(.CLK(CLK), .D(PD367), .LFSR(R367), .S(P367),.INIT(1'b0));
DEC2STCH D2S368(.CLK(CLK), .D(PD368), .LFSR(R368), .S(P368),.INIT(1'b0));
DEC2STCH D2S369(.CLK(CLK), .D(PD369), .LFSR(R369), .S(P369),.INIT(1'b0));
DEC2STCH D2S370(.CLK(CLK), .D(PD370), .LFSR(R370), .S(P370),.INIT(1'b0));
DEC2STCH D2S371(.CLK(CLK), .D(PD371), .LFSR(R371), .S(P371),.INIT(1'b0));
DEC2STCH D2S372(.CLK(CLK), .D(PD372), .LFSR(R372), .S(P372),.INIT(1'b0));
DEC2STCH D2S373(.CLK(CLK), .D(PD373), .LFSR(R373), .S(P373),.INIT(1'b0));
DEC2STCH D2S374(.CLK(CLK), .D(PD374), .LFSR(R374), .S(P374),.INIT(1'b0));
DEC2STCH D2S375(.CLK(CLK), .D(PD375), .LFSR(R375), .S(P375),.INIT(1'b0));
DEC2STCH D2S376(.CLK(CLK), .D(PD376), .LFSR(R376), .S(P376),.INIT(1'b0));
DEC2STCH D2S377(.CLK(CLK), .D(PD377), .LFSR(R377), .S(P377),.INIT(1'b0));
DEC2STCH D2S378(.CLK(CLK), .D(PD378), .LFSR(R378), .S(P378),.INIT(1'b0));
DEC2STCH D2S379(.CLK(CLK), .D(PD379), .LFSR(R379), .S(P379),.INIT(1'b0));
DEC2STCH D2S380(.CLK(CLK), .D(PD380), .LFSR(R380), .S(P380),.INIT(1'b0));
DEC2STCH D2S381(.CLK(CLK), .D(PD381), .LFSR(R381), .S(P381),.INIT(1'b0));
DEC2STCH D2S382(.CLK(CLK), .D(PD382), .LFSR(R382), .S(P382),.INIT(1'b0));
DEC2STCH D2S383(.CLK(CLK), .D(PD383), .LFSR(R383), .S(P383),.INIT(1'b0));
DEC2STCH D2S384(.CLK(CLK), .D(PD384), .LFSR(R384), .S(P384),.INIT(1'b0));
DEC2STCH D2S385(.CLK(CLK), .D(PD385), .LFSR(R385), .S(P385),.INIT(1'b0));
DEC2STCH D2S386(.CLK(CLK), .D(PD386), .LFSR(R386), .S(P386),.INIT(1'b0));
DEC2STCH D2S387(.CLK(CLK), .D(PD387), .LFSR(R387), .S(P387),.INIT(1'b0));
DEC2STCH D2S388(.CLK(CLK), .D(PD388), .LFSR(R388), .S(P388),.INIT(1'b0));
DEC2STCH D2S389(.CLK(CLK), .D(PD389), .LFSR(R389), .S(P389),.INIT(1'b0));
DEC2STCH D2S390(.CLK(CLK), .D(PD390), .LFSR(R390), .S(P390),.INIT(1'b0));
DEC2STCH D2S391(.CLK(CLK), .D(PD391), .LFSR(R391), .S(P391),.INIT(1'b0));
DEC2STCH D2S392(.CLK(CLK), .D(PD392), .LFSR(R392), .S(P392),.INIT(1'b0));
DEC2STCH D2S393(.CLK(CLK), .D(PD393), .LFSR(R393), .S(P393),.INIT(1'b0));
DEC2STCH D2S394(.CLK(CLK), .D(PD394), .LFSR(R394), .S(P394),.INIT(1'b0));
DEC2STCH D2S395(.CLK(CLK), .D(PD395), .LFSR(R395), .S(P395),.INIT(1'b0));
DEC2STCH D2S396(.CLK(CLK), .D(PD396), .LFSR(R396), .S(P396),.INIT(1'b0));
DEC2STCH D2S397(.CLK(CLK), .D(PD397), .LFSR(R397), .S(P397),.INIT(1'b0));
DEC2STCH D2S398(.CLK(CLK), .D(PD398), .LFSR(R398), .S(P398),.INIT(1'b0));
DEC2STCH D2S399(.CLK(CLK), .D(PD399), .LFSR(R399), .S(P399),.INIT(1'b0));
DEC2STCH D2S400(.CLK(CLK), .D(PD400), .LFSR(R400), .S(P400),.INIT(1'b0));
DEC2STCH D2S401(.CLK(CLK), .D(PD401), .LFSR(R401), .S(P401),.INIT(1'b0));
DEC2STCH D2S402(.CLK(CLK), .D(PD402), .LFSR(R402), .S(P402),.INIT(1'b0));
DEC2STCH D2S403(.CLK(CLK), .D(PD403), .LFSR(R403), .S(P403),.INIT(1'b0));
DEC2STCH D2S404(.CLK(CLK), .D(PD404), .LFSR(R404), .S(P404),.INIT(1'b0));
DEC2STCH D2S405(.CLK(CLK), .D(PD405), .LFSR(R405), .S(P405),.INIT(1'b0));
DEC2STCH D2S406(.CLK(CLK), .D(PD406), .LFSR(R406), .S(P406),.INIT(1'b0));
DEC2STCH D2S407(.CLK(CLK), .D(PD407), .LFSR(R407), .S(P407),.INIT(1'b0));
DEC2STCH D2S408(.CLK(CLK), .D(PD408), .LFSR(R408), .S(P408),.INIT(1'b0));
DEC2STCH D2S409(.CLK(CLK), .D(PD409), .LFSR(R409), .S(P409),.INIT(1'b0));
DEC2STCH D2S410(.CLK(CLK), .D(PD410), .LFSR(R410), .S(P410),.INIT(1'b0));
DEC2STCH D2S411(.CLK(CLK), .D(PD411), .LFSR(R411), .S(P411),.INIT(1'b0));
DEC2STCH D2S412(.CLK(CLK), .D(PD412), .LFSR(R412), .S(P412),.INIT(1'b0));
DEC2STCH D2S413(.CLK(CLK), .D(PD413), .LFSR(R413), .S(P413),.INIT(1'b0));
DEC2STCH D2S414(.CLK(CLK), .D(PD414), .LFSR(R414), .S(P414),.INIT(1'b0));
DEC2STCH D2S415(.CLK(CLK), .D(PD415), .LFSR(R415), .S(P415),.INIT(1'b0));
DEC2STCH D2S416(.CLK(CLK), .D(PD416), .LFSR(R416), .S(P416),.INIT(1'b0));
DEC2STCH D2S417(.CLK(CLK), .D(PD417), .LFSR(R417), .S(P417),.INIT(1'b0));
DEC2STCH D2S418(.CLK(CLK), .D(PD418), .LFSR(R418), .S(P418),.INIT(1'b0));
DEC2STCH D2S419(.CLK(CLK), .D(PD419), .LFSR(R419), .S(P419),.INIT(1'b0));
DEC2STCH D2S420(.CLK(CLK), .D(PD420), .LFSR(R420), .S(P420),.INIT(1'b0));
DEC2STCH D2S421(.CLK(CLK), .D(PD421), .LFSR(R421), .S(P421),.INIT(1'b0));
DEC2STCH D2S422(.CLK(CLK), .D(PD422), .LFSR(R422), .S(P422),.INIT(1'b0));
DEC2STCH D2S423(.CLK(CLK), .D(PD423), .LFSR(R423), .S(P423),.INIT(1'b0));
DEC2STCH D2S424(.CLK(CLK), .D(PD424), .LFSR(R424), .S(P424),.INIT(1'b0));
DEC2STCH D2S425(.CLK(CLK), .D(PD425), .LFSR(R425), .S(P425),.INIT(1'b0));
DEC2STCH D2S426(.CLK(CLK), .D(PD426), .LFSR(R426), .S(P426),.INIT(1'b0));
DEC2STCH D2S427(.CLK(CLK), .D(PD427), .LFSR(R427), .S(P427),.INIT(1'b0));
DEC2STCH D2S428(.CLK(CLK), .D(PD428), .LFSR(R428), .S(P428),.INIT(1'b0));
DEC2STCH D2S429(.CLK(CLK), .D(PD429), .LFSR(R429), .S(P429),.INIT(1'b0));
DEC2STCH D2S430(.CLK(CLK), .D(PD430), .LFSR(R430), .S(P430),.INIT(1'b0));
DEC2STCH D2S431(.CLK(CLK), .D(PD431), .LFSR(R431), .S(P431),.INIT(1'b0));
DEC2STCH D2S432(.CLK(CLK), .D(PD432), .LFSR(R432), .S(P432),.INIT(1'b0));
DEC2STCH D2S433(.CLK(CLK), .D(PD433), .LFSR(R433), .S(P433),.INIT(1'b0));
DEC2STCH D2S434(.CLK(CLK), .D(PD434), .LFSR(R434), .S(P434),.INIT(1'b0));
DEC2STCH D2S435(.CLK(CLK), .D(PD435), .LFSR(R435), .S(P435),.INIT(1'b0));
DEC2STCH D2S436(.CLK(CLK), .D(PD436), .LFSR(R436), .S(P436),.INIT(1'b0));
DEC2STCH D2S437(.CLK(CLK), .D(PD437), .LFSR(R437), .S(P437),.INIT(1'b0));
DEC2STCH D2S438(.CLK(CLK), .D(PD438), .LFSR(R438), .S(P438),.INIT(1'b0));
DEC2STCH D2S439(.CLK(CLK), .D(PD439), .LFSR(R439), .S(P439),.INIT(1'b0));
DEC2STCH D2S440(.CLK(CLK), .D(PD440), .LFSR(R440), .S(P440),.INIT(1'b0));
DEC2STCH D2S441(.CLK(CLK), .D(PD441), .LFSR(R441), .S(P441),.INIT(1'b0));
DEC2STCH D2S442(.CLK(CLK), .D(PD442), .LFSR(R442), .S(P442),.INIT(1'b0));
DEC2STCH D2S443(.CLK(CLK), .D(PD443), .LFSR(R443), .S(P443),.INIT(1'b0));
DEC2STCH D2S444(.CLK(CLK), .D(PD444), .LFSR(R444), .S(P444),.INIT(1'b0));
DEC2STCH D2S445(.CLK(CLK), .D(PD445), .LFSR(R445), .S(P445),.INIT(1'b0));
DEC2STCH D2S446(.CLK(CLK), .D(PD446), .LFSR(R446), .S(P446),.INIT(1'b0));
DEC2STCH D2S447(.CLK(CLK), .D(PD447), .LFSR(R447), .S(P447),.INIT(1'b0));
DEC2STCH D2S448(.CLK(CLK), .D(PD448), .LFSR(R448), .S(P448),.INIT(1'b0));
DEC2STCH D2S449(.CLK(CLK), .D(PD449), .LFSR(R449), .S(P449),.INIT(1'b0));
DEC2STCH D2S450(.CLK(CLK), .D(PD450), .LFSR(R450), .S(P450),.INIT(1'b0));
DEC2STCH D2S451(.CLK(CLK), .D(PD451), .LFSR(R451), .S(P451),.INIT(1'b0));
DEC2STCH D2S452(.CLK(CLK), .D(PD452), .LFSR(R452), .S(P452),.INIT(1'b0));
DEC2STCH D2S453(.CLK(CLK), .D(PD453), .LFSR(R453), .S(P453),.INIT(1'b0));
DEC2STCH D2S454(.CLK(CLK), .D(PD454), .LFSR(R454), .S(P454),.INIT(1'b0));
DEC2STCH D2S455(.CLK(CLK), .D(PD455), .LFSR(R455), .S(P455),.INIT(1'b0));
DEC2STCH D2S456(.CLK(CLK), .D(PD456), .LFSR(R456), .S(P456),.INIT(1'b0));

// Long D2S Conversion:

DEC2STCH D2S_long0(.CLK(CLK), .D(PD_long0), .LFSR(R_long0), .S(P_long0),.INIT(1'b0));
DEC2STCH D2S_long1(.CLK(CLK), .D(PD_long1), .LFSR(R_long1), .S(P_long1),.INIT(1'b0));
DEC2STCH D2S_long2(.CLK(CLK), .D(PD_long2), .LFSR(R_long2), .S(P_long2),.INIT(1'b0));
DEC2STCH D2S_long3(.CLK(CLK), .D(PD_long3), .LFSR(R_long3), .S(P_long3),.INIT(1'b0));
DEC2STCH D2S_long4(.CLK(CLK), .D(PD_long4), .LFSR(R_long4), .S(P_long4),.INIT(1'b0));
DEC2STCH D2S_long5(.CLK(CLK), .D(PD_long5), .LFSR(R_long5), .S(P_long5),.INIT(1'b0));
DEC2STCH D2S_long6(.CLK(CLK), .D(PD_long6), .LFSR(R_long6), .S(P_long6),.INIT(1'b0));
DEC2STCH D2S_long7(.CLK(CLK), .D(PD_long7), .LFSR(R_long7), .S(P_long7),.INIT(1'b0));
DEC2STCH D2S_long8(.CLK(CLK), .D(PD_long8), .LFSR(R_long8), .S(P_long8),.INIT(1'b0));
DEC2STCH D2S_long9(.CLK(CLK), .D(PD_long9), .LFSR(R_long9), .S(P_long9),.INIT(1'b0));
DEC2STCH D2S_long10(.CLK(CLK), .D(PD_long10), .LFSR(R_long10), .S(P_long10),.INIT(1'b0));
DEC2STCH D2S_long11(.CLK(CLK), .D(PD_long11), .LFSR(R_long11), .S(P_long11),.INIT(1'b0));
DEC2STCH D2S_long12(.CLK(CLK), .D(PD_long12), .LFSR(R_long12), .S(P_long12),.INIT(1'b0));
DEC2STCH D2S_long13(.CLK(CLK), .D(PD_long13), .LFSR(R_long13), .S(P_long13),.INIT(1'b0));
DEC2STCH D2S_long14(.CLK(CLK), .D(PD_long14), .LFSR(R_long14), .S(P_long14),.INIT(1'b0));
defparam D2S_long0.ND = DP_out;
defparam D2S_long1.ND = DP_out;
defparam D2S_long2.ND = DP_out;
defparam D2S_long3.ND = DP_out;
defparam D2S_long4.ND = DP_out;
defparam D2S_long5.ND = DP_out;
defparam D2S_long6.ND = DP_out;
defparam D2S_long7.ND = DP_out;
defparam D2S_long8.ND = DP_out;
defparam D2S_long9.ND = DP_out;
defparam D2S_long10.ND = DP_out;
defparam D2S_long11.ND = DP_out;
defparam D2S_long12.ND = DP_out;
defparam D2S_long13.ND = DP_out;
defparam D2S_long14.ND = DP_out;

endmodule